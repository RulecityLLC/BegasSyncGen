--------------------------------------------------------------------------------
-- Company: 	RuleCity LLC
-- Engineer:	Matt Ownby

-- NOTE: run simulator to at least 5 uS to cover all test cases.

--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY outputGenTest IS
END outputGenTest;
 
ARCHITECTURE behavior OF outputGenTest IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT outputGen
    PORT(
         clock14_3 : IN  std_logic;
			reset_prime : IN std_logic;
         is_top_field : OUT  boolean;
			subcarrier_out : out  STD_LOGIC;
         sgblk_prime : OUT  std_logic;
         hsync2_prime : OUT  std_logic;
			csync_prime : OUT  std_logic;
         vsync2_prime : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clock14_3 : std_logic := '0';
	signal reset_prime : std_logic := '1';

 	--Outputs
   signal is_top_field : boolean;
	signal subcarrier_out : std_logic;
   signal sgblk_prime : std_logic;
   signal hsync2_prime : std_logic;
	signal csync_prime : std_logic;
   signal vsync2_prime : std_logic;

   -- Clock period definitions
   constant clock14_3_period : time := 10 ps;	-- smaller is more convenient

BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: outputGen PORT MAP (
          clock14_3 => clock14_3,
			 reset_prime => reset_prime,
          is_top_field => is_top_field,
			 subcarrier_out => subcarrier_out,
          sgblk_prime => sgblk_prime,
          hsync2_prime => hsync2_prime,
			 csync_prime => csync_prime,
          vsync2_prime => vsync2_prime
        );

   -- Clock process definitions
   clock14_3_process :process
   begin
		-- easier to debug if we start at 1
		clock14_3 <= '1';
		wait for clock14_3_period/2;
		clock14_3 <= '0';
		wait for clock14_3_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		

		-- sub carrier test
		wait for clock14_3_period;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime (SC test)" severity failure;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime (SC test)" severity failure;
		assert (subcarrier_out = '1') report "Unexpected value for subcarrier (SC test)" severity failure;

		wait for clock14_3_period;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime (SC test)" severity failure;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime (SC test)" severity failure;
		assert (subcarrier_out = '1') report "Unexpected value for subcarrier (SC test)" severity failure;

		wait for clock14_3_period;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime (SC test)" severity failure;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime (SC test)" severity failure;
		assert (subcarrier_out = '0') report "Unexpected value for subcarrier (SC test)" severity failure;

		wait for clock14_3_period;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime (SC test)" severity failure;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime (SC test)" severity failure;
		assert (subcarrier_out = '0') report "Unexpected value for subcarrier (SC test)" severity failure;
		
		-- test reset

		wait for clock14_3_period * 8296;	-- somewhat arbitrary, puts us in area where hsync and vsync are both disabled
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime" severity failure;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime" severity failure;

		-- reset should move us back to 0 after a single clock cycle
		reset_prime <= '0';
		wait for clock14_3_period;
		reset_prime <= '1';

		-- *** AUTO GENERATED CODE FOLLOWS ***


		--next cycle transition
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 0" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 0" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 0" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 21" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 21" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 21" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 22" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 53" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 53" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 53" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 53" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 54" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 95" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 95" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 95" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 95" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 96" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 476" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 476" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 476" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 476" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 477" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 508" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 508" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 508" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 508" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 509" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 909" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 909" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 909" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 931" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 931" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 931" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 931" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 932" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 963" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 963" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 963" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 963" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 964" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 1005" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 1005" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 1005" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 1005" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 1006" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 1386" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 1386" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 1386" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 1386" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 1387" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 1418" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 1418" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 1418" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 1418" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 1419" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 1819" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 1819" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 1819" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 1819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 1820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 1841" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 1841" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 1841" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 1841" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 1842" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 1873" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 1873" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 1873" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 1873" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 1874" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 1915" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 1915" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 1915" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 1915" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 1916" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 2296" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 2296" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 2296" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 2296" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 2297" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 2328" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 2328" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 2328" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 2328" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 2329" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 2729" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 2729" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 2729" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 2729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 2730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 2751" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 2751" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 2751" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 2751" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 2752" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 73);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 2825" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 2825" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 2825" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 2825" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 2826" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 312);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 3138" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 3138" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 3138" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 3138" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 3139" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 3206" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 3206" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 3206" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 3206" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 3207" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 386);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 3593" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 3593" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 3593" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 3593" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 3594" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 45);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 3639" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 3639" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 3639" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 3639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 3640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 3661" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 3661" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 3661" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 3661" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 3662" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 73);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 3735" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 3735" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 3735" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 3735" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 3736" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 312);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 4048" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 4048" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 4048" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 4048" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 4049" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 4116" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 4116" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 4116" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 4116" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 4117" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 386);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 4503" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 4503" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 4503" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 4503" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 4504" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 45);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 4549" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 4549" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 4549" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 4549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 4550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 4571" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 4571" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 4571" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 4571" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 4572" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 73);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 4645" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 4645" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 4645" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 4645" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 4646" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 312);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 4958" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 4958" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 4958" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 4958" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 4959" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 5026" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 5026" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 5026" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 5026" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 5027" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 386);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 5413" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 5413" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 5413" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 5413" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 5414" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 45);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 5459" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 5459" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 5459" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 5459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 5460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 5481" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 5481" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 5481" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 5481" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 5482" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 5513" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 5513" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 5513" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 5513" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 5514" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 5555" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 5555" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 5555" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 5555" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 5556" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 5936" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 5936" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 5936" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 5936" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 5937" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 5968" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 5968" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 5968" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 5968" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 5969" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 6369" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 6369" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 6369" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 6369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 6370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 6391" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 6391" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 6391" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 6391" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 6392" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 6423" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 6423" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 6423" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 6423" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 6424" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 6465" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 6465" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 6465" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 6465" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 6466" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 6846" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 6846" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 6846" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 6846" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 6847" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 6878" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 6878" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 6878" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 6878" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 6879" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 7279" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 7279" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 7279" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 7279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 7280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 7301" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 7301" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 7301" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 7301" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 7302" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 7333" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 7333" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 7333" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 7333" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 7334" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 7375" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 7375" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 7375" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 7375" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 7376" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 7756" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 7756" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 7756" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 7756" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 7757" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 7788" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 7788" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 7788" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 7788" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 7789" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 8189" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 8189" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 8189" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 8189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 8190" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 8190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 8211" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 8211" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 8211" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 8211" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 8212" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 8279" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 8279" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 8279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 8279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 8280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 8285" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 8285" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 8285" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 8285" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 8286" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 9099" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 9099" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 9099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 9099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 9100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 9121" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 9121" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 9121" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 9121" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 9122" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 9189" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 9189" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 9189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 9189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 9190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 9195" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 9195" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 9195" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 9195" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 9196" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 10009" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 10009" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 10009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 10009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 10010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 10031" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 10031" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 10031" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 10031" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 10032" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 10099" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 10099" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 10099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 10099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 10100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 10105" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 10105" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 10105" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 10105" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 10106" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 10919" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 10919" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 10919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 10919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 10920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 10941" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 10941" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 10941" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 10941" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 10942" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 11009" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 11009" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 11009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 11009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 11010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 11015" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 11015" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 11015" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 11015" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 11016" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 11829" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 11829" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 11829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 11829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 11830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 11851" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 11851" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 11851" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 11851" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 11852" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 11919" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 11919" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 11919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 11919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 11920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 11925" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 11925" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 11925" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 11925" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 11926" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 12739" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 12739" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 12739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 12739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 12740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 12761" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 12761" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 12761" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 12761" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 12762" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 12829" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 12829" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 12829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 12829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 12830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 12835" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 12835" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 12835" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 12835" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 12836" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 13649" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 13649" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 13649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 13649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 13650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 13671" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 13671" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 13671" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 13671" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 13672" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 13739" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 13739" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 13739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 13739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 13740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 13745" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 13745" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 13745" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 13745" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 13746" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 14559" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 14559" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 14559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 14559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 14560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 14581" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 14581" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 14581" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 14581" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 14582" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 14649" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 14649" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 14649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 14649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 14650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 14655" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 14655" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 14655" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 14655" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 14656" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 15469" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 15469" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 15469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 15469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 15470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 15491" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 15491" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 15491" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 15491" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 15492" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 15559" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 15559" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 15559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 15559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 15560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 15565" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 15565" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 15565" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 15565" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 15566" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 16379" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 16379" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 16379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 16379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 16380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 16401" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 16401" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 16401" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 16401" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 16402" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 16469" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 16469" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 16469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 16469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 16470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 16475" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 16475" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 16475" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 16475" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 16476" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 17289" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 17289" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 17289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 17289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 17290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 17311" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 17311" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 17311" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 17311" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 17312" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 17379" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 17379" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 17379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 17379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 17380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 17385" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 17385" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 17385" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 17385" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 17386" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 18199" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 18199" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 18199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 18199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 18200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 18221" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 18221" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 18221" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 18221" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 18222" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 18289" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 18289" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 18289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 18289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 18290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 18295" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 18295" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 18295" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 18295" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 18296" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 18353" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 18353" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 18353" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 18353" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 18354" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 19109" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 19109" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 19109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 19109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 19110" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 19110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 19131" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 19131" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 19131" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 19131" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 19132" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 19199" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 19199" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 19199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 19199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 19200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 19205" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 19205" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 19205" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 19205" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 19206" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 19263" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 19263" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 19263" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 19263" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 19264" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 20019" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 20019" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 20019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 20019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 20020" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 20020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 20041" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 20041" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 20041" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 20041" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 20042" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 20109" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 20109" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 20109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 20109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 20110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 20115" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 20115" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 20115" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 20115" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 20116" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 20173" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 20173" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 20173" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 20173" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 20174" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 20929" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 20929" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 20929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 20929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 20930" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 20930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 20951" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 20951" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 20951" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 20951" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 20952" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 21019" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 21019" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 21019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 21019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 21020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 21025" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 21025" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 21025" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 21025" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 21026" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 21083" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 21083" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 21083" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 21083" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 21084" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 21839" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 21839" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 21839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 21839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 21840" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 21840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 21861" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 21861" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 21861" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 21861" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 21862" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 21929" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 21929" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 21929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 21929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 21930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 21935" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 21935" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 21935" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 21935" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 21936" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 21993" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 21993" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 21993" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 21993" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 21994" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 22749" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 22749" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 22749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 22749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 22750" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 22750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 22771" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 22771" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 22771" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 22771" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 22772" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 22839" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 22839" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 22839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 22839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 22840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 22845" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 22845" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 22845" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 22845" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 22846" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 22903" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 22903" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 22903" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 22903" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 22904" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 23659" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 23659" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 23659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 23659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 23660" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 23660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 23681" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 23681" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 23681" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 23681" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 23682" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 23749" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 23749" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 23749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 23749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 23750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 23755" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 23755" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 23755" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 23755" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 23756" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 23813" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 23813" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 23813" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 23813" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 23814" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 24569" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 24569" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 24569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 24569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 24570" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 24570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 24591" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 24591" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 24591" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 24591" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 24592" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 24659" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 24659" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 24659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 24659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 24660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 24665" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 24665" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 24665" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 24665" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 24666" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 24723" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 24723" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 24723" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 24723" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 24724" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 25479" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 25479" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 25479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 25479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 25480" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 25480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 25501" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 25501" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 25501" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 25501" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 25502" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 25569" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 25569" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 25569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 25569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 25570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 25575" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 25575" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 25575" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 25575" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 25576" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 25633" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 25633" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 25633" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 25633" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 25634" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 26389" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 26389" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 26389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 26389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 26390" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 26390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 26411" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 26411" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 26411" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 26411" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 26412" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 26479" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 26479" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 26479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 26479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 26480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 26485" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 26485" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 26485" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 26485" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 26486" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 26543" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 26543" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 26543" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 26543" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 26544" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 27299" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 27299" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 27299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 27299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 27300" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 27300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 27321" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 27321" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 27321" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 27321" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 27322" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 27389" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 27389" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 27389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 27389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 27390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 27395" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 27395" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 27395" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 27395" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 27396" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 27453" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 27453" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 27453" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 27453" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 27454" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 28209" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 28209" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 28209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 28209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 28210" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 28210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 28231" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 28231" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 28231" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 28231" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 28232" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 28299" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 28299" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 28299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 28299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 28300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 28305" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 28305" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 28305" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 28305" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 28306" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 28363" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 28363" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 28363" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 28363" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 28364" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 29119" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 29119" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 29119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 29119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 29120" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 29120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 29141" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 29141" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 29141" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 29141" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 29142" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 29209" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 29209" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 29209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 29209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 29210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 29215" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 29215" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 29215" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 29215" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 29216" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 29273" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 29273" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 29273" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 29273" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 29274" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 30029" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 30029" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 30029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 30029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 30030" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 30030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 30051" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 30051" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 30051" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 30051" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 30052" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 30119" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 30119" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 30119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 30119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 30120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 30125" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 30125" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 30125" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 30125" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 30126" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 30183" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 30183" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 30183" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 30183" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 30184" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 30939" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 30939" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 30939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 30939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 30940" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 30940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 30961" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 30961" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 30961" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 30961" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 30962" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 31029" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 31029" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 31029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 31029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 31030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 31035" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 31035" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 31035" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 31035" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 31036" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 31093" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 31093" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 31093" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 31093" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 31094" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 31849" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 31849" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 31849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 31849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 31850" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 31850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 31871" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 31871" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 31871" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 31871" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 31872" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 31939" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 31939" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 31939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 31939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 31940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 31945" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 31945" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 31945" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 31945" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 31946" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 32003" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 32003" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 32003" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 32003" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 32004" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 32759" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 32759" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 32759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 32759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 32760" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 32760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 32781" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 32781" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 32781" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 32781" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 32782" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 32849" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 32849" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 32849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 32849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 32850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 32855" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 32855" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 32855" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 32855" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 32856" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 32913" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 32913" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 32913" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 32913" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 32914" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 33669" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 33669" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 33669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 33669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 33670" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 33670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 33691" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 33691" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 33691" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 33691" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 33692" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 33759" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 33759" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 33759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 33759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 33760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 33765" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 33765" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 33765" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 33765" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 33766" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 33823" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 33823" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 33823" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 33823" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 33824" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 34579" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 34579" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 34579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 34579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 34580" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 34580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 34601" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 34601" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 34601" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 34601" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 34602" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 34669" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 34669" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 34669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 34669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 34670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 34675" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 34675" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 34675" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 34675" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 34676" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 34733" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 34733" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 34733" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 34733" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 34734" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 35489" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 35489" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 35489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 35489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 35490" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 35490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 35511" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 35511" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 35511" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 35511" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 35512" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 35579" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 35579" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 35579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 35579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 35580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 35585" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 35585" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 35585" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 35585" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 35586" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 35643" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 35643" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 35643" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 35643" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 35644" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 36399" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 36399" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 36399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 36399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 36400" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 36400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 36421" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 36421" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 36421" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 36421" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 36422" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 36489" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 36489" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 36489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 36489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 36490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 36495" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 36495" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 36495" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 36495" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 36496" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 36553" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 36553" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 36553" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 36553" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 36554" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 37309" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 37309" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 37309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 37309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 37310" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 37310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 37331" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 37331" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 37331" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 37331" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 37332" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 37399" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 37399" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 37399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 37399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 37400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 37405" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 37405" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 37405" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 37405" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 37406" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 37463" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 37463" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 37463" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 37463" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 37464" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 38219" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 38219" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 38219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 38219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 38220" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 38220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 38241" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 38241" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 38241" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 38241" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 38242" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 38309" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 38309" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 38309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 38309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 38310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 38315" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 38315" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 38315" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 38315" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 38316" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 38373" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 38373" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 38373" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 38373" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 38374" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 39129" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 39129" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 39129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 39129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 39130" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 39130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 39151" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 39151" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 39151" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 39151" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 39152" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 39219" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 39219" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 39219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 39219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 39220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 39225" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 39225" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 39225" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 39225" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 39226" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 39283" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 39283" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 39283" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 39283" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 39284" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 40039" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 40039" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 40039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 40039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 40040" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 40040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 40061" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 40061" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 40061" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 40061" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 40062" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 40129" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 40129" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 40129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 40129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 40130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 40135" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 40135" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 40135" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 40135" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 40136" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 40193" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 40193" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 40193" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 40193" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 40194" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 40949" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 40949" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 40949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 40949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 40950" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 40950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 40971" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 40971" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 40971" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 40971" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 40972" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 41039" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 41039" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 41039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 41039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 41040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 41045" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 41045" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 41045" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 41045" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 41046" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 41103" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 41103" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 41103" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 41103" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 41104" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 41859" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 41859" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 41859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 41859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 41860" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 41860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 41881" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 41881" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 41881" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 41881" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 41882" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 41949" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 41949" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 41949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 41949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 41950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 41955" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 41955" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 41955" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 41955" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 41956" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 42013" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 42013" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 42013" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 42013" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 42014" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 42769" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 42769" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 42769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 42769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 42770" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 42770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 42791" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 42791" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 42791" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 42791" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 42792" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 42859" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 42859" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 42859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 42859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 42860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 42865" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 42865" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 42865" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 42865" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 42866" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 42923" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 42923" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 42923" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 42923" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 42924" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 43679" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 43679" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 43679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 43679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 43680" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 43680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 43701" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 43701" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 43701" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 43701" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 43702" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 43769" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 43769" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 43769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 43769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 43770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 43775" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 43775" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 43775" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 43775" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 43776" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 43833" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 43833" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 43833" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 43833" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 43834" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 44589" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 44589" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 44589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 44589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 44590" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 44590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 44611" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 44611" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 44611" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 44611" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 44612" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 44679" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 44679" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 44679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 44679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 44680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 44685" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 44685" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 44685" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 44685" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 44686" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 44743" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 44743" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 44743" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 44743" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 44744" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 45499" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 45499" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 45499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 45499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 45500" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 45500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 45521" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 45521" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 45521" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 45521" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 45522" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 45589" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 45589" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 45589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 45589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 45590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 45595" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 45595" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 45595" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 45595" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 45596" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 45653" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 45653" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 45653" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 45653" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 45654" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 46409" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 46409" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 46409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 46409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 46410" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 46410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 46431" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 46431" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 46431" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 46431" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 46432" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 46499" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 46499" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 46499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 46499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 46500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 46505" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 46505" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 46505" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 46505" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 46506" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 46563" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 46563" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 46563" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 46563" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 46564" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 47319" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 47319" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 47319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 47319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 47320" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 47320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 47341" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 47341" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 47341" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 47341" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 47342" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 47409" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 47409" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 47409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 47409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 47410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 47415" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 47415" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 47415" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 47415" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 47416" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 47473" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 47473" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 47473" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 47473" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 47474" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 48229" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 48229" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 48229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 48229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 48230" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 48230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 48251" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 48251" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 48251" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 48251" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 48252" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 48319" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 48319" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 48319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 48319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 48320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 48325" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 48325" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 48325" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 48325" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 48326" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 48383" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 48383" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 48383" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 48383" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 48384" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 49139" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 49139" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 49139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 49139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 49140" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 49140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 49161" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 49161" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 49161" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 49161" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 49162" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 49229" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 49229" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 49229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 49229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 49230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 49235" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 49235" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 49235" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 49235" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 49236" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 49293" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 49293" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 49293" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 49293" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 49294" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 50049" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 50049" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 50049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 50049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 50050" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 50050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 50071" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 50071" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 50071" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 50071" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 50072" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 50139" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 50139" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 50139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 50139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 50140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 50145" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 50145" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 50145" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 50145" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 50146" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 50203" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 50203" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 50203" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 50203" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 50204" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 50959" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 50959" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 50959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 50959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 50960" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 50960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 50981" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 50981" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 50981" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 50981" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 50982" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 51049" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 51049" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 51049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 51049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 51050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 51055" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 51055" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 51055" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 51055" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 51056" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 51113" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 51113" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 51113" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 51113" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 51114" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 51869" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 51869" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 51869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 51869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 51870" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 51870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 51891" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 51891" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 51891" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 51891" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 51892" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 51959" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 51959" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 51959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 51959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 51960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 51965" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 51965" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 51965" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 51965" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 51966" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 52023" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 52023" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 52023" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 52023" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 52024" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 52779" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 52779" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 52779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 52779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 52780" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 52780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 52801" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 52801" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 52801" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 52801" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 52802" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 52869" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 52869" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 52869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 52869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 52870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 52875" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 52875" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 52875" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 52875" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 52876" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 52933" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 52933" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 52933" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 52933" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 52934" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 53689" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 53689" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 53689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 53689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 53690" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 53690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 53711" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 53711" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 53711" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 53711" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 53712" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 53779" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 53779" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 53779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 53779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 53780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 53785" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 53785" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 53785" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 53785" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 53786" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 53843" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 53843" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 53843" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 53843" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 53844" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 54599" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 54599" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 54599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 54599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 54600" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 54600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 54621" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 54621" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 54621" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 54621" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 54622" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 54689" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 54689" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 54689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 54689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 54690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 54695" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 54695" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 54695" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 54695" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 54696" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 54753" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 54753" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 54753" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 54753" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 54754" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 55509" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 55509" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 55509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 55509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 55510" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 55510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 55531" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 55531" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 55531" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 55531" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 55532" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 55599" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 55599" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 55599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 55599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 55600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 55605" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 55605" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 55605" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 55605" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 55606" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 55663" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 55663" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 55663" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 55663" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 55664" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 56419" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 56419" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 56419" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 56419" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 56420" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 56420" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 56441" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 56441" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 56441" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 56441" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 56442" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 56509" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 56509" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 56509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 56509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 56510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 56515" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 56515" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 56515" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 56515" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 56516" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 56573" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 56573" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 56573" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 56573" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 56574" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 57329" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 57329" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 57329" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 57329" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 57330" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 57330" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 57351" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 57351" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 57351" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 57351" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 57352" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 57419" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 57419" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 57419" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 57419" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 57420" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 57425" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 57425" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 57425" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 57425" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 57426" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 57483" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 57483" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 57483" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 57483" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 57484" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 58239" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 58239" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 58239" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 58239" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 58240" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 58240" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 58261" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 58261" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 58261" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 58261" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 58262" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 58329" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 58329" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 58329" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 58329" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 58330" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 58335" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 58335" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 58335" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 58335" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 58336" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 58393" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 58393" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 58393" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 58393" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 58394" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 59149" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 59149" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 59149" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 59149" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 59150" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 59150" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 59171" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 59171" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 59171" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 59171" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 59172" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 59239" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 59239" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 59239" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 59239" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 59240" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 59245" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 59245" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 59245" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 59245" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 59246" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 59303" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 59303" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 59303" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 59303" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 59304" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 60059" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 60059" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 60059" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 60059" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 60060" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 60060" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 60081" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 60081" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 60081" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 60081" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 60082" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 60149" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 60149" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 60149" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 60149" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 60150" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 60155" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 60155" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 60155" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 60155" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 60156" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 60213" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 60213" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 60213" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 60213" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 60214" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 60969" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 60969" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 60969" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 60969" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 60970" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 60970" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 60991" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 60991" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 60991" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 60991" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 60992" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 61059" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 61059" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 61059" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 61059" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 61060" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 61065" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 61065" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 61065" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 61065" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 61066" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 61123" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 61123" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 61123" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 61123" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 61124" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 61879" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 61879" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 61879" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 61879" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 61880" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 61880" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 61901" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 61901" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 61901" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 61901" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 61902" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 61969" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 61969" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 61969" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 61969" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 61970" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 61975" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 61975" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 61975" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 61975" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 61976" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 62033" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 62033" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 62033" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 62033" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 62034" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 62789" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 62789" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 62789" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 62789" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 62790" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 62790" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 62811" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 62811" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 62811" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 62811" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 62812" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 62879" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 62879" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 62879" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 62879" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 62880" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 62885" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 62885" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 62885" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 62885" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 62886" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 62943" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 62943" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 62943" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 62943" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 62944" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 63699" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 63699" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 63699" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 63699" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 63700" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 63700" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 63721" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 63721" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 63721" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 63721" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 63722" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 63789" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 63789" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 63789" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 63789" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 63790" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 63795" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 63795" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 63795" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 63795" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 63796" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 63853" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 63853" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 63853" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 63853" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 63854" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 64609" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 64609" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 64609" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 64609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 64610" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 64610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 64631" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 64631" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 64631" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 64631" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 64632" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 64699" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 64699" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 64699" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 64699" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 64700" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 64705" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 64705" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 64705" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 64705" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 64706" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 64763" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 64763" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 64763" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 64763" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 64764" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 65519" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 65519" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 65519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 65519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 65520" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 65520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 65541" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 65541" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 65541" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 65541" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 65542" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 65609" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 65609" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 65609" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 65609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 65610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 65615" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 65615" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 65615" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 65615" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 65616" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 65673" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 65673" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 65673" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 65673" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 65674" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 66429" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 66429" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 66429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 66429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 66430" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 66430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 66451" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 66451" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 66451" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 66451" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 66452" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 66519" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 66519" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 66519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 66519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 66520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 66525" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 66525" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 66525" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 66525" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 66526" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 66583" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 66583" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 66583" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 66583" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 66584" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 67339" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 67339" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 67339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 67339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 67340" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 67340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 67361" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 67361" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 67361" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 67361" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 67362" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 67429" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 67429" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 67429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 67429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 67430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 67435" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 67435" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 67435" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 67435" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 67436" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 67493" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 67493" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 67493" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 67493" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 67494" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 68249" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 68249" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 68249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 68249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 68250" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 68250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 68271" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 68271" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 68271" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 68271" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 68272" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 68339" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 68339" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 68339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 68339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 68340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 68345" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 68345" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 68345" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 68345" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 68346" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 68403" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 68403" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 68403" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 68403" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 68404" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 69159" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 69159" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 69159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 69159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 69160" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 69160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 69181" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 69181" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 69181" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 69181" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 69182" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 69249" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 69249" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 69249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 69249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 69250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 69255" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 69255" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 69255" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 69255" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 69256" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 69313" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 69313" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 69313" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 69313" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 69314" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 70069" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 70069" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 70069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 70069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 70070" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 70070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 70091" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 70091" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 70091" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 70091" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 70092" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 70159" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 70159" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 70159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 70159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 70160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 70165" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 70165" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 70165" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 70165" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 70166" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 70223" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 70223" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 70223" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 70223" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 70224" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 70979" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 70979" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 70979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 70979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 70980" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 70980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 71001" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 71001" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 71001" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 71001" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 71002" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 71069" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 71069" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 71069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 71069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 71070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 71075" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 71075" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 71075" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 71075" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 71076" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 71133" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 71133" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 71133" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 71133" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 71134" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 71889" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 71889" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 71889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 71889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 71890" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 71890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 71911" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 71911" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 71911" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 71911" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 71912" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 71979" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 71979" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 71979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 71979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 71980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 71985" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 71985" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 71985" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 71985" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 71986" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 72043" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 72043" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 72043" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 72043" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 72044" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 72799" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 72799" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 72799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 72799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 72800" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 72800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 72821" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 72821" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 72821" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 72821" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 72822" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 72889" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 72889" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 72889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 72889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 72890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 72895" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 72895" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 72895" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 72895" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 72896" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 72953" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 72953" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 72953" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 72953" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 72954" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 73709" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 73709" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 73709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 73709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 73710" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 73710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 73731" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 73731" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 73731" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 73731" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 73732" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 73799" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 73799" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 73799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 73799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 73800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 73805" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 73805" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 73805" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 73805" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 73806" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 73863" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 73863" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 73863" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 73863" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 73864" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 74619" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 74619" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 74619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 74619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 74620" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 74620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 74641" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 74641" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 74641" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 74641" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 74642" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 74709" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 74709" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 74709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 74709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 74710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 74715" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 74715" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 74715" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 74715" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 74716" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 74773" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 74773" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 74773" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 74773" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 74774" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 75529" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 75529" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 75529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 75529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 75530" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 75530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 75551" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 75551" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 75551" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 75551" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 75552" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 75619" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 75619" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 75619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 75619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 75620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 75625" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 75625" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 75625" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 75625" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 75626" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 75683" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 75683" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 75683" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 75683" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 75684" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 76439" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 76439" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 76439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 76439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 76440" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 76440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 76461" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 76461" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 76461" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 76461" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 76462" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 76529" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 76529" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 76529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 76529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 76530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 76535" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 76535" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 76535" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 76535" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 76536" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 76593" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 76593" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 76593" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 76593" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 76594" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 77349" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 77349" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 77349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 77349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 77350" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 77350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 77371" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 77371" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 77371" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 77371" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 77372" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 77439" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 77439" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 77439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 77439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 77440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 77445" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 77445" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 77445" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 77445" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 77446" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 77503" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 77503" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 77503" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 77503" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 77504" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 78259" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 78259" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 78259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 78259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 78260" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 78260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 78281" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 78281" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 78281" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 78281" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 78282" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 78349" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 78349" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 78349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 78349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 78350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 78355" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 78355" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 78355" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 78355" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 78356" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 78413" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 78413" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 78413" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 78413" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 78414" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 79169" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 79169" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 79169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 79169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 79170" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 79170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 79191" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 79191" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 79191" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 79191" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 79192" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 79259" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 79259" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 79259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 79259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 79260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 79265" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 79265" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 79265" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 79265" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 79266" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 79323" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 79323" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 79323" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 79323" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 79324" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 80079" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 80079" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 80079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 80079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 80080" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 80080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 80101" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 80101" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 80101" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 80101" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 80102" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 80169" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 80169" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 80169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 80169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 80170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 80175" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 80175" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 80175" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 80175" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 80176" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 80233" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 80233" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 80233" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 80233" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 80234" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 80989" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 80989" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 80989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 80989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 80990" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 80990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 81011" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 81011" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 81011" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 81011" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 81012" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 81079" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 81079" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 81079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 81079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 81080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 81085" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 81085" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 81085" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 81085" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 81086" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 81143" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 81143" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 81143" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 81143" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 81144" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 81899" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 81899" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 81899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 81899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 81900" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 81900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 81921" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 81921" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 81921" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 81921" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 81922" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 81989" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 81989" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 81989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 81989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 81990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 81995" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 81995" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 81995" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 81995" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 81996" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 82053" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 82053" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 82053" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 82053" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 82054" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 82809" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 82809" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 82809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 82809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 82810" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 82810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 82831" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 82831" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 82831" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 82831" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 82832" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 82899" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 82899" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 82899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 82899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 82900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 82905" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 82905" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 82905" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 82905" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 82906" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 82963" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 82963" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 82963" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 82963" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 82964" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 83719" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 83719" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 83719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 83719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 83720" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 83720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 83741" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 83741" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 83741" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 83741" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 83742" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 83809" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 83809" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 83809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 83809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 83810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 83815" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 83815" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 83815" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 83815" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 83816" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 83873" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 83873" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 83873" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 83873" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 83874" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 84629" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 84629" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 84629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 84629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 84630" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 84630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 84651" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 84651" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 84651" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 84651" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 84652" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 84719" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 84719" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 84719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 84719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 84720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 84725" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 84725" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 84725" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 84725" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 84726" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 84783" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 84783" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 84783" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 84783" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 84784" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 85539" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 85539" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 85539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 85539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 85540" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 85540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 85561" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 85561" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 85561" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 85561" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 85562" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 85629" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 85629" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 85629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 85629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 85630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 85635" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 85635" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 85635" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 85635" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 85636" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 85693" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 85693" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 85693" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 85693" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 85694" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 86449" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 86449" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 86449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 86449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 86450" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 86450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 86471" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 86471" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 86471" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 86471" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 86472" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 86539" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 86539" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 86539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 86539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 86540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 86545" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 86545" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 86545" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 86545" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 86546" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 86603" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 86603" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 86603" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 86603" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 86604" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 87359" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 87359" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 87359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 87359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 87360" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 87360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 87381" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 87381" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 87381" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 87381" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 87382" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 87449" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 87449" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 87449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 87449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 87450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 87455" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 87455" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 87455" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 87455" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 87456" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 87513" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 87513" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 87513" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 87513" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 87514" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 88269" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 88269" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 88269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 88269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 88270" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 88270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 88291" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 88291" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 88291" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 88291" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 88292" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 88359" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 88359" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 88359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 88359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 88360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 88365" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 88365" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 88365" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 88365" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 88366" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 88423" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 88423" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 88423" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 88423" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 88424" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 89179" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 89179" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 89179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 89179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 89180" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 89180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 89201" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 89201" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 89201" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 89201" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 89202" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 89269" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 89269" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 89269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 89269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 89270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 89275" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 89275" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 89275" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 89275" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 89276" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 89333" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 89333" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 89333" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 89333" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 89334" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 90089" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 90089" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 90089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 90089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 90090" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 90090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 90111" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 90111" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 90111" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 90111" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 90112" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 90179" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 90179" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 90179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 90179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 90180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 90185" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 90185" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 90185" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 90185" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 90186" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 90243" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 90243" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 90243" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 90243" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 90244" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 90999" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 90999" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 90999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 90999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 91000" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 91000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 91021" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 91021" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 91021" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 91021" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 91022" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 91089" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 91089" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 91089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 91089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 91090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 91095" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 91095" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 91095" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 91095" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 91096" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 91153" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 91153" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 91153" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 91153" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 91154" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 91909" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 91909" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 91909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 91909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 91910" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 91910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 91931" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 91931" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 91931" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 91931" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 91932" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 91999" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 91999" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 91999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 91999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 92000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 92005" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 92005" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 92005" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 92005" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 92006" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 92063" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 92063" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 92063" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 92063" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 92064" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 92819" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 92819" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 92819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 92819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 92820" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 92820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 92841" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 92841" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 92841" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 92841" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 92842" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 92909" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 92909" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 92909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 92909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 92910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 92915" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 92915" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 92915" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 92915" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 92916" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 92973" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 92973" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 92973" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 92973" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 92974" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 93729" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 93729" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 93729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 93729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 93730" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 93730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 93751" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 93751" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 93751" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 93751" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 93752" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 93819" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 93819" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 93819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 93819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 93820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 93825" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 93825" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 93825" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 93825" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 93826" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 93883" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 93883" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 93883" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 93883" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 93884" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 94639" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 94639" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 94639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 94639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 94640" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 94640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 94661" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 94661" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 94661" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 94661" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 94662" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 94729" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 94729" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 94729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 94729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 94730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 94735" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 94735" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 94735" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 94735" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 94736" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 94793" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 94793" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 94793" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 94793" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 94794" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 95549" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 95549" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 95549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 95549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 95550" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 95550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 95571" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 95571" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 95571" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 95571" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 95572" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 95639" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 95639" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 95639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 95639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 95640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 95645" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 95645" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 95645" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 95645" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 95646" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 95703" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 95703" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 95703" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 95703" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 95704" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 96459" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 96459" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 96459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 96459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 96460" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 96460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 96481" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 96481" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 96481" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 96481" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 96482" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 96549" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 96549" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 96549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 96549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 96550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 96555" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 96555" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 96555" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 96555" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 96556" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 96613" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 96613" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 96613" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 96613" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 96614" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 97369" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 97369" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 97369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 97369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 97370" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 97370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 97391" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 97391" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 97391" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 97391" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 97392" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 97459" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 97459" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 97459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 97459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 97460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 97465" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 97465" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 97465" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 97465" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 97466" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 97523" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 97523" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 97523" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 97523" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 97524" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 98279" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 98279" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 98279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 98279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 98280" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 98280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 98301" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 98301" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 98301" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 98301" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 98302" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 98369" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 98369" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 98369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 98369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 98370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 98375" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 98375" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 98375" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 98375" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 98376" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 98433" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 98433" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 98433" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 98433" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 98434" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 99189" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 99189" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 99189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 99189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 99190" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 99190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 99211" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 99211" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 99211" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 99211" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 99212" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 99279" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 99279" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 99279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 99279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 99280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 99285" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 99285" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 99285" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 99285" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 99286" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 99343" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 99343" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 99343" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 99343" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 99344" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 100099" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 100099" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 100099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 100099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 100100" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 100100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 100121" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 100121" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 100121" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 100121" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 100122" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 100189" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 100189" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 100189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 100189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 100190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 100195" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 100195" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 100195" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 100195" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 100196" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 100253" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 100253" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 100253" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 100253" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 100254" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 101009" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 101009" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 101009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 101009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 101010" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 101010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 101031" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 101031" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 101031" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 101031" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 101032" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 101099" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 101099" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 101099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 101099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 101100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 101105" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 101105" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 101105" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 101105" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 101106" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 101163" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 101163" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 101163" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 101163" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 101164" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 101919" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 101919" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 101919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 101919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 101920" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 101920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 101941" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 101941" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 101941" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 101941" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 101942" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 102009" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 102009" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 102009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 102009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 102010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 102015" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 102015" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 102015" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 102015" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 102016" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 102073" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 102073" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 102073" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 102073" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 102074" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 102829" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 102829" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 102829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 102829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 102830" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 102830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 102851" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 102851" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 102851" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 102851" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 102852" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 102919" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 102919" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 102919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 102919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 102920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 102925" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 102925" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 102925" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 102925" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 102926" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 102983" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 102983" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 102983" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 102983" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 102984" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 103739" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 103739" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 103739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 103739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 103740" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 103740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 103761" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 103761" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 103761" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 103761" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 103762" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 103829" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 103829" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 103829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 103829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 103830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 103835" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 103835" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 103835" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 103835" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 103836" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 103893" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 103893" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 103893" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 103893" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 103894" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 104649" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 104649" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 104649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 104649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 104650" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 104650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 104671" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 104671" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 104671" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 104671" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 104672" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 104739" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 104739" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 104739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 104739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 104740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 104745" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 104745" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 104745" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 104745" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 104746" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 104803" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 104803" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 104803" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 104803" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 104804" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 105559" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 105559" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 105559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 105559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 105560" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 105560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 105581" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 105581" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 105581" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 105581" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 105582" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 105649" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 105649" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 105649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 105649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 105650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 105655" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 105655" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 105655" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 105655" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 105656" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 105713" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 105713" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 105713" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 105713" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 105714" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 106469" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 106469" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 106469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 106469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 106470" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 106470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 106491" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 106491" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 106491" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 106491" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 106492" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 106559" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 106559" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 106559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 106559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 106560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 106565" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 106565" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 106565" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 106565" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 106566" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 106623" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 106623" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 106623" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 106623" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 106624" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 107379" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 107379" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 107379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 107379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 107380" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 107380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 107401" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 107401" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 107401" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 107401" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 107402" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 107469" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 107469" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 107469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 107469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 107470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 107475" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 107475" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 107475" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 107475" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 107476" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 107533" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 107533" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 107533" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 107533" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 107534" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 108289" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 108289" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 108289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 108289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 108290" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 108290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 108311" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 108311" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 108311" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 108311" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 108312" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 108379" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 108379" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 108379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 108379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 108380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 108385" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 108385" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 108385" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 108385" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 108386" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 108443" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 108443" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 108443" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 108443" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 108444" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 109199" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 109199" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 109199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 109199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 109200" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 109200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 109221" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 109221" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 109221" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 109221" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 109222" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 109289" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 109289" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 109289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 109289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 109290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 109295" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 109295" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 109295" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 109295" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 109296" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 109353" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 109353" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 109353" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 109353" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 109354" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 110109" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 110109" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 110109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 110109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 110110" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 110110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 110131" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 110131" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 110131" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 110131" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 110132" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 110199" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 110199" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 110199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 110199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 110200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 110205" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 110205" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 110205" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 110205" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 110206" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 110263" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 110263" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 110263" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 110263" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 110264" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 111019" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 111019" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 111019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 111019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 111020" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 111020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 111041" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 111041" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 111041" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 111041" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 111042" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 111109" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 111109" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 111109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 111109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 111110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 111115" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 111115" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 111115" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 111115" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 111116" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 111173" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 111173" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 111173" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 111173" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 111174" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 111929" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 111929" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 111929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 111929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 111930" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 111930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 111951" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 111951" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 111951" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 111951" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 111952" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 112019" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 112019" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 112019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 112019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 112020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 112025" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 112025" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 112025" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 112025" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 112026" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 112083" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 112083" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 112083" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 112083" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 112084" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 112839" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 112839" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 112839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 112839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 112840" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 112840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 112861" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 112861" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 112861" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 112861" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 112862" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 112929" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 112929" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 112929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 112929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 112930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 112935" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 112935" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 112935" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 112935" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 112936" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 112993" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 112993" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 112993" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 112993" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 112994" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 113749" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 113749" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 113749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 113749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 113750" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 113750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 113771" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 113771" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 113771" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 113771" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 113772" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 113839" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 113839" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 113839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 113839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 113840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 113845" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 113845" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 113845" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 113845" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 113846" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 113903" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 113903" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 113903" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 113903" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 113904" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 114659" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 114659" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 114659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 114659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 114660" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 114660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 114681" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 114681" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 114681" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 114681" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 114682" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 114749" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 114749" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 114749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 114749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 114750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 114755" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 114755" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 114755" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 114755" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 114756" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 114813" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 114813" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 114813" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 114813" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 114814" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 115569" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 115569" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 115569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 115569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 115570" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 115570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 115591" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 115591" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 115591" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 115591" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 115592" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 115659" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 115659" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 115659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 115659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 115660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 115665" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 115665" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 115665" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 115665" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 115666" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 115723" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 115723" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 115723" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 115723" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 115724" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 116479" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 116479" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 116479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 116479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 116480" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 116480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 116501" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 116501" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 116501" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 116501" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 116502" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 116569" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 116569" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 116569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 116569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 116570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 116575" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 116575" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 116575" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 116575" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 116576" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 116633" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 116633" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 116633" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 116633" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 116634" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 117389" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 117389" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 117389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 117389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 117390" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 117390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 117411" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 117411" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 117411" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 117411" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 117412" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 117479" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 117479" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 117479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 117479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 117480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 117485" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 117485" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 117485" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 117485" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 117486" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 117543" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 117543" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 117543" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 117543" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 117544" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 118299" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 118299" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 118299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 118299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 118300" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 118300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 118321" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 118321" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 118321" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 118321" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 118322" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 118389" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 118389" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 118389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 118389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 118390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 118395" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 118395" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 118395" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 118395" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 118396" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 118453" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 118453" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 118453" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 118453" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 118454" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 119209" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 119209" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 119209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 119209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 119210" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 119210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 119231" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 119231" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 119231" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 119231" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 119232" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 119299" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 119299" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 119299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 119299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 119300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 119305" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 119305" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 119305" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 119305" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 119306" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 119363" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 119363" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 119363" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 119363" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 119364" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 120119" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 120119" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 120119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 120119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 120120" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 120120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 120141" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 120141" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 120141" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 120141" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 120142" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 120209" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 120209" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 120209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 120209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 120210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 120215" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 120215" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 120215" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 120215" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 120216" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 120273" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 120273" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 120273" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 120273" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 120274" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 121029" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 121029" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 121029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 121029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 121030" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 121030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 121051" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 121051" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 121051" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 121051" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 121052" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 121119" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 121119" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 121119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 121119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 121120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 121125" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 121125" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 121125" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 121125" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 121126" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 121183" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 121183" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 121183" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 121183" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 121184" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 121939" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 121939" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 121939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 121939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 121940" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 121940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 121961" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 121961" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 121961" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 121961" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 121962" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 122029" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 122029" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 122029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 122029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 122030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 122035" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 122035" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 122035" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 122035" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 122036" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 122093" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 122093" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 122093" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 122093" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 122094" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 122849" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 122849" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 122849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 122849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 122850" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 122850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 122871" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 122871" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 122871" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 122871" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 122872" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 122939" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 122939" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 122939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 122939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 122940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 122945" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 122945" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 122945" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 122945" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 122946" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 123003" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 123003" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 123003" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 123003" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 123004" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 123759" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 123759" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 123759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 123759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 123760" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 123760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 123781" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 123781" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 123781" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 123781" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 123782" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 123849" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 123849" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 123849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 123849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 123850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 123855" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 123855" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 123855" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 123855" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 123856" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 123913" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 123913" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 123913" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 123913" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 123914" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 124669" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 124669" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 124669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 124669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 124670" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 124670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 124691" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 124691" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 124691" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 124691" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 124692" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 124759" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 124759" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 124759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 124759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 124760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 124765" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 124765" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 124765" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 124765" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 124766" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 124823" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 124823" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 124823" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 124823" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 124824" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 125579" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 125579" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 125579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 125579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 125580" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 125580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 125601" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 125601" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 125601" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 125601" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 125602" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 125669" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 125669" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 125669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 125669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 125670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 125675" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 125675" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 125675" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 125675" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 125676" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 125733" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 125733" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 125733" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 125733" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 125734" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 126489" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 126489" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 126489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 126489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 126490" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 126490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 126511" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 126511" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 126511" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 126511" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 126512" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 126579" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 126579" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 126579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 126579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 126580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 126585" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 126585" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 126585" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 126585" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 126586" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 126643" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 126643" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 126643" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 126643" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 126644" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 127399" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 127399" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 127399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 127399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 127400" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 127400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 127421" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 127421" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 127421" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 127421" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 127422" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 127489" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 127489" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 127489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 127489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 127490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 127495" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 127495" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 127495" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 127495" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 127496" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 127553" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 127553" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 127553" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 127553" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 127554" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 128309" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 128309" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 128309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 128309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 128310" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 128310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 128331" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 128331" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 128331" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 128331" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 128332" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 128399" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 128399" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 128399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 128399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 128400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 128405" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 128405" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 128405" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 128405" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 128406" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 128463" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 128463" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 128463" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 128463" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 128464" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 129219" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 129219" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 129219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 129219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 129220" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 129220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 129241" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 129241" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 129241" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 129241" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 129242" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 129309" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 129309" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 129309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 129309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 129310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 129315" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 129315" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 129315" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 129315" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 129316" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 129373" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 129373" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 129373" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 129373" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 129374" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 130129" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 130129" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 130129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 130129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 130130" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 130130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 130151" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 130151" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 130151" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 130151" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 130152" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 130219" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 130219" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 130219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 130219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 130220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 130225" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 130225" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 130225" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 130225" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 130226" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 130283" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 130283" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 130283" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 130283" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 130284" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 131039" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 131039" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 131039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 131039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 131040" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 131040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 131061" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 131061" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 131061" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 131061" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 131062" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 131129" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 131129" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 131129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 131129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 131130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 131135" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 131135" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 131135" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 131135" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 131136" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 131193" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 131193" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 131193" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 131193" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 131194" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 131949" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 131949" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 131949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 131949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 131950" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 131950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 131971" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 131971" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 131971" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 131971" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 131972" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 132039" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 132039" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 132039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 132039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 132040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 132045" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 132045" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 132045" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 132045" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 132046" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 132103" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 132103" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 132103" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 132103" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 132104" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 132859" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 132859" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 132859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 132859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 132860" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 132860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 132881" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 132881" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 132881" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 132881" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 132882" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 132949" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 132949" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 132949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 132949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 132950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 132955" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 132955" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 132955" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 132955" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 132956" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 133013" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 133013" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 133013" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 133013" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 133014" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 133769" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 133769" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 133769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 133769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 133770" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 133770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 133791" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 133791" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 133791" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 133791" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 133792" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 133859" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 133859" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 133859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 133859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 133860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 133865" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 133865" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 133865" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 133865" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 133866" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 133923" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 133923" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 133923" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 133923" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 133924" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 134679" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 134679" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 134679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 134679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 134680" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 134680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 134701" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 134701" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 134701" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 134701" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 134702" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 134769" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 134769" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 134769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 134769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 134770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 134775" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 134775" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 134775" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 134775" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 134776" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 134833" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 134833" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 134833" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 134833" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 134834" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 135589" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 135589" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 135589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 135589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 135590" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 135590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 135611" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 135611" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 135611" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 135611" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 135612" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 135679" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 135679" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 135679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 135679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 135680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 135685" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 135685" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 135685" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 135685" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 135686" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 135743" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 135743" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 135743" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 135743" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 135744" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 136499" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 136499" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 136499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 136499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 136500" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 136500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 136521" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 136521" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 136521" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 136521" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 136522" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 136589" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 136589" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 136589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 136589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 136590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 136595" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 136595" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 136595" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 136595" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 136596" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 136653" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 136653" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 136653" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 136653" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 136654" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 137409" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 137409" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 137409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 137409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 137410" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 137410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 137431" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 137431" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 137431" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 137431" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 137432" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 137499" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 137499" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 137499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 137499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 137500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 137505" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 137505" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 137505" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 137505" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 137506" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 137563" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 137563" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 137563" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 137563" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 137564" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 138319" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 138319" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 138319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 138319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 138320" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 138320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 138341" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 138341" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 138341" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 138341" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 138342" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 138409" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 138409" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 138409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 138409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 138410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 138415" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 138415" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 138415" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 138415" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 138416" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 138473" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 138473" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 138473" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 138473" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 138474" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 139229" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 139229" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 139229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 139229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 139230" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 139230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 139251" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 139251" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 139251" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 139251" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 139252" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 139319" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 139319" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 139319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 139319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 139320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 139325" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 139325" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 139325" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 139325" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 139326" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 139383" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 139383" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 139383" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 139383" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 139384" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 140139" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 140139" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 140139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 140139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 140140" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 140140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 140161" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 140161" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 140161" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 140161" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 140162" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 140229" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 140229" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 140229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 140229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 140230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 140235" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 140235" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 140235" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 140235" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 140236" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 140293" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 140293" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 140293" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 140293" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 140294" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 141049" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 141049" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 141049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 141049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 141050" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 141050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 141071" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 141071" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 141071" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 141071" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 141072" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 141139" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 141139" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 141139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 141139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 141140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 141145" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 141145" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 141145" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 141145" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 141146" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 141203" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 141203" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 141203" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 141203" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 141204" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 141959" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 141959" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 141959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 141959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 141960" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 141960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 141981" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 141981" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 141981" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 141981" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 141982" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 142049" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 142049" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 142049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 142049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 142050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 142055" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 142055" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 142055" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 142055" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 142056" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 142113" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 142113" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 142113" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 142113" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 142114" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 142869" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 142869" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 142869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 142869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 142870" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 142870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 142891" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 142891" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 142891" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 142891" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 142892" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 142959" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 142959" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 142959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 142959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 142960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 142965" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 142965" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 142965" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 142965" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 142966" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 143023" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 143023" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 143023" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 143023" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 143024" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 143779" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 143779" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 143779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 143779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 143780" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 143780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 143801" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 143801" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 143801" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 143801" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 143802" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 143869" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 143869" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 143869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 143869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 143870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 143875" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 143875" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 143875" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 143875" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 143876" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 143933" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 143933" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 143933" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 143933" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 143934" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 144689" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 144689" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 144689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 144689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 144690" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 144690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 144711" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 144711" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 144711" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 144711" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 144712" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 144779" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 144779" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 144779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 144779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 144780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 144785" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 144785" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 144785" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 144785" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 144786" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 144843" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 144843" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 144843" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 144843" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 144844" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 145599" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 145599" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 145599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 145599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 145600" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 145600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 145621" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 145621" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 145621" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 145621" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 145622" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 145689" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 145689" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 145689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 145689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 145690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 145695" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 145695" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 145695" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 145695" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 145696" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 145753" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 145753" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 145753" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 145753" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 145754" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 146509" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 146509" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 146509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 146509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 146510" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 146510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 146531" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 146531" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 146531" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 146531" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 146532" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 146599" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 146599" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 146599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 146599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 146600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 146605" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 146605" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 146605" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 146605" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 146606" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 146663" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 146663" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 146663" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 146663" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 146664" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 147419" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 147419" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 147419" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 147419" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 147420" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 147420" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 147441" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 147441" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 147441" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 147441" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 147442" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 147509" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 147509" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 147509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 147509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 147510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 147515" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 147515" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 147515" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 147515" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 147516" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 147573" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 147573" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 147573" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 147573" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 147574" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 148329" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 148329" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 148329" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 148329" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 148330" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 148330" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 148351" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 148351" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 148351" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 148351" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 148352" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 148419" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 148419" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 148419" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 148419" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 148420" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 148425" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 148425" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 148425" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 148425" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 148426" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 148483" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 148483" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 148483" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 148483" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 148484" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 149239" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 149239" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 149239" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 149239" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 149240" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 149240" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 149261" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 149261" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 149261" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 149261" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 149262" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 149329" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 149329" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 149329" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 149329" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 149330" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 149335" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 149335" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 149335" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 149335" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 149336" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 149393" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 149393" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 149393" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 149393" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 149394" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 150149" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 150149" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 150149" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 150149" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 150150" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 150150" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 150171" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 150171" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 150171" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 150171" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 150172" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 150239" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 150239" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 150239" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 150239" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 150240" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 150245" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 150245" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 150245" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 150245" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 150246" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 150303" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 150303" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 150303" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 150303" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 150304" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 151059" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 151059" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 151059" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 151059" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 151060" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 151060" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 151081" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 151081" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 151081" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 151081" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 151082" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 151149" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 151149" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 151149" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 151149" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 151150" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 151155" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 151155" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 151155" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 151155" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 151156" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 151213" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 151213" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 151213" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 151213" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 151214" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 151969" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 151969" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 151969" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 151969" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 151970" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 151970" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 151991" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 151991" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 151991" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 151991" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 151992" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 152059" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 152059" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 152059" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 152059" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 152060" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 152065" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 152065" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 152065" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 152065" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 152066" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 152123" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 152123" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 152123" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 152123" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 152124" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 152879" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 152879" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 152879" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 152879" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 152880" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 152880" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 152901" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 152901" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 152901" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 152901" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 152902" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 152969" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 152969" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 152969" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 152969" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 152970" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 152975" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 152975" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 152975" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 152975" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 152976" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 153033" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 153033" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 153033" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 153033" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 153034" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 153789" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 153789" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 153789" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 153789" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 153790" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 153790" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 153811" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 153811" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 153811" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 153811" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 153812" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 153879" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 153879" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 153879" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 153879" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 153880" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 153885" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 153885" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 153885" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 153885" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 153886" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 153943" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 153943" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 153943" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 153943" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 153944" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 154699" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 154699" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 154699" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 154699" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 154700" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 154700" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 154721" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 154721" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 154721" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 154721" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 154722" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 154789" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 154789" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 154789" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 154789" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 154790" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 154795" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 154795" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 154795" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 154795" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 154796" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 154853" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 154853" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 154853" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 154853" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 154854" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 155609" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 155609" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 155609" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 155609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 155610" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 155610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 155631" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 155631" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 155631" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 155631" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 155632" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 155699" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 155699" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 155699" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 155699" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 155700" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 155705" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 155705" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 155705" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 155705" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 155706" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 155763" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 155763" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 155763" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 155763" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 155764" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 156519" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 156519" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 156519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 156519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 156520" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 156520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 156541" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 156541" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 156541" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 156541" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 156542" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 156609" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 156609" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 156609" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 156609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 156610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 156615" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 156615" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 156615" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 156615" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 156616" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 156673" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 156673" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 156673" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 156673" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 156674" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 157429" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 157429" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 157429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 157429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 157430" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 157430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 157451" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 157451" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 157451" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 157451" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 157452" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 157519" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 157519" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 157519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 157519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 157520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 157525" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 157525" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 157525" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 157525" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 157526" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 157583" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 157583" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 157583" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 157583" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 157584" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 158339" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 158339" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 158339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 158339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 158340" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 158340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 158361" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 158361" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 158361" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 158361" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 158362" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 158429" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 158429" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 158429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 158429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 158430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 158435" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 158435" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 158435" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 158435" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 158436" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 158493" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 158493" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 158493" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 158493" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 158494" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 159249" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 159249" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 159249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 159249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 159250" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 159250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 159271" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 159271" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 159271" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 159271" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 159272" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 159339" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 159339" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 159339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 159339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 159340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 159345" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 159345" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 159345" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 159345" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 159346" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 159403" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 159403" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 159403" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 159403" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 159404" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 160159" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 160159" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 160159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 160159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 160160" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 160160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 160181" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 160181" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 160181" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 160181" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 160182" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 160249" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 160249" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 160249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 160249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 160250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 160255" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 160255" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 160255" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 160255" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 160256" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 160313" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 160313" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 160313" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 160313" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 160314" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 161069" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 161069" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 161069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 161069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 161070" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 161070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 161091" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 161091" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 161091" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 161091" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 161092" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 161159" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 161159" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 161159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 161159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 161160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 161165" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 161165" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 161165" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 161165" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 161166" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 161223" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 161223" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 161223" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 161223" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 161224" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 161979" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 161979" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 161979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 161979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 161980" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 161980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 162001" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 162001" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 162001" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 162001" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 162002" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 162069" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 162069" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 162069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 162069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 162070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 162075" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 162075" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 162075" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 162075" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 162076" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 162133" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 162133" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 162133" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 162133" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 162134" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 162889" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 162889" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 162889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 162889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 162890" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 162890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 162911" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 162911" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 162911" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 162911" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 162912" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 162979" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 162979" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 162979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 162979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 162980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 162985" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 162985" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 162985" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 162985" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 162986" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 163043" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 163043" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 163043" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 163043" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 163044" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 163799" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 163799" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 163799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 163799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 163800" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 163800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 163821" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 163821" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 163821" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 163821" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 163822" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 163889" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 163889" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 163889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 163889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 163890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 163895" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 163895" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 163895" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 163895" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 163896" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 163953" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 163953" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 163953" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 163953" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 163954" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 164709" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 164709" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 164709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 164709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 164710" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 164710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 164731" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 164731" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 164731" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 164731" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 164732" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 164799" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 164799" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 164799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 164799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 164800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 164805" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 164805" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 164805" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 164805" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 164806" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 164863" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 164863" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 164863" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 164863" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 164864" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 165619" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 165619" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 165619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 165619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 165620" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 165620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 165641" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 165641" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 165641" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 165641" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 165642" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 165709" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 165709" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 165709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 165709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 165710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 165715" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 165715" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 165715" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 165715" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 165716" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 165773" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 165773" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 165773" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 165773" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 165774" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 166529" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 166529" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 166529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 166529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 166530" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 166530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 166551" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 166551" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 166551" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 166551" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 166552" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 166619" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 166619" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 166619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 166619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 166620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 166625" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 166625" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 166625" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 166625" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 166626" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 166683" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 166683" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 166683" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 166683" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 166684" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 167439" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 167439" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 167439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 167439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 167440" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 167440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 167461" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 167461" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 167461" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 167461" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 167462" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 167529" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 167529" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 167529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 167529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 167530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 167535" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 167535" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 167535" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 167535" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 167536" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 167593" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 167593" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 167593" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 167593" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 167594" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 168349" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 168349" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 168349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 168349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 168350" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 168350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 168371" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 168371" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 168371" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 168371" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 168372" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 168439" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 168439" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 168439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 168439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 168440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 168445" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 168445" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 168445" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 168445" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 168446" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 168503" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 168503" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 168503" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 168503" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 168504" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 169259" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 169259" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 169259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 169259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 169260" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 169260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 169281" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 169281" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 169281" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 169281" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 169282" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 169349" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 169349" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 169349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 169349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 169350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 169355" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 169355" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 169355" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 169355" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 169356" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 169413" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 169413" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 169413" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 169413" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 169414" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 170169" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 170169" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 170169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 170169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 170170" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 170170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 170191" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 170191" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 170191" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 170191" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 170192" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 170259" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 170259" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 170259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 170259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 170260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 170265" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 170265" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 170265" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 170265" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 170266" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 170323" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 170323" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 170323" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 170323" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 170324" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 171079" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 171079" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 171079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 171079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 171080" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 171080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 171101" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 171101" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 171101" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 171101" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 171102" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 171169" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 171169" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 171169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 171169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 171170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 171175" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 171175" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 171175" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 171175" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 171176" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 171233" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 171233" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 171233" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 171233" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 171234" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 171989" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 171989" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 171989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 171989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 171990" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 171990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 172011" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 172011" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 172011" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 172011" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 172012" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 172079" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 172079" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 172079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 172079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 172080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 172085" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 172085" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 172085" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 172085" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 172086" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 172143" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 172143" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 172143" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 172143" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 172144" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 172899" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 172899" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 172899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 172899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 172900" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 172900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 172921" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 172921" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 172921" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 172921" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 172922" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 172989" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 172989" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 172989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 172989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 172990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 172995" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 172995" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 172995" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 172995" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 172996" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 173053" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 173053" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 173053" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 173053" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 173054" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 173809" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 173809" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 173809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 173809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 173810" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 173810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 173831" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 173831" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 173831" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 173831" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 173832" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 173899" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 173899" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 173899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 173899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 173900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 173905" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 173905" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 173905" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 173905" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 173906" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 173963" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 173963" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 173963" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 173963" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 173964" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 174719" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 174719" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 174719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 174719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 174720" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 174720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 174741" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 174741" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 174741" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 174741" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 174742" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 174809" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 174809" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 174809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 174809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 174810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 174815" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 174815" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 174815" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 174815" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 174816" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 174873" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 174873" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 174873" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 174873" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 174874" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 175629" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 175629" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 175629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 175629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 175630" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 175630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 175651" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 175651" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 175651" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 175651" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 175652" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 175719" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 175719" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 175719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 175719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 175720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 175725" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 175725" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 175725" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 175725" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 175726" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 175783" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 175783" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 175783" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 175783" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 175784" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 176539" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 176539" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 176539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 176539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 176540" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 176540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 176561" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 176561" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 176561" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 176561" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 176562" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 176629" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 176629" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 176629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 176629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 176630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 176635" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 176635" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 176635" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 176635" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 176636" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 176693" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 176693" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 176693" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 176693" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 176694" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 177449" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 177449" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 177449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 177449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 177450" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 177450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 177471" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 177471" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 177471" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 177471" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 177472" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 177539" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 177539" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 177539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 177539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 177540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 177545" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 177545" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 177545" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 177545" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 177546" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 177603" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 177603" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 177603" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 177603" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 177604" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 178359" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 178359" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 178359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 178359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 178360" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 178360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 178381" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 178381" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 178381" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 178381" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 178382" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 178449" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 178449" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 178449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 178449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 178450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 178455" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 178455" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 178455" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 178455" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 178456" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 178513" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 178513" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 178513" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 178513" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 178514" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 179269" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 179269" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 179269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 179269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 179270" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 179270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 179291" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 179291" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 179291" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 179291" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 179292" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 179359" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 179359" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 179359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 179359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 179360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 179365" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 179365" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 179365" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 179365" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 179366" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 179423" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 179423" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 179423" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 179423" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 179424" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 180179" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 180179" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 180179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 180179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 180180" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 180180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 180201" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 180201" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 180201" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 180201" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 180202" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 180269" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 180269" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 180269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 180269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 180270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 180275" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 180275" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 180275" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 180275" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 180276" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 180333" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 180333" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 180333" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 180333" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 180334" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 181089" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 181089" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 181089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 181089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 181090" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 181090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 181111" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 181111" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 181111" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 181111" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 181112" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 181179" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 181179" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 181179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 181179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 181180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 181185" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 181185" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 181185" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 181185" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 181186" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 181243" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 181243" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 181243" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 181243" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 181244" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 181999" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 181999" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 181999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 181999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 182000" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 182000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 182021" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 182021" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 182021" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 182021" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 182022" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 182089" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 182089" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 182089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 182089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 182090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 182095" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 182095" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 182095" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 182095" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 182096" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 182153" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 182153" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 182153" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 182153" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 182154" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 182909" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 182909" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 182909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 182909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 182910" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 182910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 182931" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 182931" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 182931" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 182931" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 182932" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 182999" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 182999" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 182999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 182999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 183000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 183005" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 183005" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 183005" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 183005" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 183006" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 183063" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 183063" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 183063" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 183063" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 183064" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 183819" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 183819" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 183819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 183819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 183820" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 183820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 183841" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 183841" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 183841" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 183841" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 183842" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 183909" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 183909" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 183909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 183909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 183910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 183915" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 183915" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 183915" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 183915" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 183916" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 183973" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 183973" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 183973" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 183973" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 183974" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 184729" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 184729" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 184729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 184729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 184730" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 184730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 184751" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 184751" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 184751" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 184751" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 184752" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 184819" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 184819" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 184819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 184819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 184820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 184825" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 184825" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 184825" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 184825" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 184826" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 184883" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 184883" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 184883" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 184883" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 184884" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 185639" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 185639" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 185639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 185639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 185640" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 185640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 185661" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 185661" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 185661" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 185661" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 185662" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 185729" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 185729" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 185729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 185729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 185730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 185735" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 185735" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 185735" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 185735" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 185736" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 185793" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 185793" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 185793" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 185793" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 185794" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 186549" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 186549" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 186549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 186549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 186550" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 186550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 186571" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 186571" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 186571" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 186571" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 186572" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 186639" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 186639" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 186639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 186639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 186640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 186645" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 186645" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 186645" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 186645" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 186646" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 186703" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 186703" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 186703" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 186703" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 186704" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 187459" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 187459" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 187459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 187459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 187460" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 187460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 187481" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 187481" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 187481" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 187481" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 187482" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 187549" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 187549" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 187549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 187549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 187550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 187555" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 187555" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 187555" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 187555" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 187556" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 187613" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 187613" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 187613" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 187613" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 187614" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 188369" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 188369" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 188369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 188369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 188370" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 188370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 188391" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 188391" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 188391" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 188391" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 188392" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 188459" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 188459" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 188459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 188459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 188460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 188465" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 188465" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 188465" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 188465" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 188466" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 188523" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 188523" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 188523" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 188523" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 188524" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 189279" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 189279" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 189279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 189279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 189280" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 189280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 189301" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 189301" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 189301" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 189301" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 189302" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 189369" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 189369" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 189369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 189369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 189370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 189375" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 189375" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 189375" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 189375" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 189376" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 189433" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 189433" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 189433" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 189433" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 189434" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 190189" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 190189" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 190189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 190189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 190190" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 190190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 190211" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 190211" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 190211" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 190211" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 190212" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 190279" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 190279" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 190279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 190279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 190280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 190285" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 190285" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 190285" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 190285" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 190286" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 190343" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 190343" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 190343" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 190343" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 190344" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 191099" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 191099" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 191099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 191099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 191100" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 191100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 191121" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 191121" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 191121" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 191121" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 191122" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 191189" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 191189" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 191189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 191189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 191190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 191195" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 191195" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 191195" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 191195" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 191196" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 191253" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 191253" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 191253" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 191253" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 191254" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 192009" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 192009" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 192009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 192009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 192010" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 192010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 192031" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 192031" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 192031" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 192031" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 192032" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 192099" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 192099" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 192099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 192099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 192100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 192105" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 192105" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 192105" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 192105" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 192106" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 192163" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 192163" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 192163" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 192163" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 192164" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 192919" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 192919" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 192919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 192919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 192920" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 192920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 192941" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 192941" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 192941" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 192941" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 192942" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 193009" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 193009" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 193009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 193009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 193010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 193015" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 193015" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 193015" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 193015" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 193016" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 193073" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 193073" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 193073" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 193073" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 193074" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 193829" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 193829" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 193829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 193829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 193830" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 193830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 193851" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 193851" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 193851" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 193851" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 193852" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 193919" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 193919" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 193919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 193919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 193920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 193925" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 193925" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 193925" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 193925" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 193926" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 193983" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 193983" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 193983" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 193983" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 193984" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 194739" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 194739" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 194739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 194739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 194740" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 194740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 194761" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 194761" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 194761" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 194761" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 194762" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 194829" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 194829" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 194829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 194829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 194830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 194835" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 194835" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 194835" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 194835" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 194836" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 194893" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 194893" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 194893" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 194893" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 194894" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 195649" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 195649" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 195649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 195649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 195650" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 195650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 195671" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 195671" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 195671" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 195671" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 195672" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 195739" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 195739" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 195739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 195739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 195740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 195745" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 195745" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 195745" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 195745" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 195746" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 195803" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 195803" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 195803" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 195803" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 195804" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 196559" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 196559" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 196559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 196559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 196560" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 196560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 196581" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 196581" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 196581" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 196581" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 196582" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 196649" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 196649" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 196649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 196649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 196650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 196655" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 196655" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 196655" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 196655" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 196656" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 196713" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 196713" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 196713" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 196713" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 196714" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 197469" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 197469" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 197469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 197469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 197470" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 197470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 197491" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 197491" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 197491" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 197491" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 197492" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 197559" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 197559" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 197559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 197559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 197560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 197565" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 197565" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 197565" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 197565" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 197566" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 197623" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 197623" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 197623" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 197623" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 197624" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 198379" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 198379" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 198379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 198379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 198380" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 198380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 198401" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 198401" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 198401" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 198401" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 198402" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 198469" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 198469" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 198469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 198469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 198470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 198475" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 198475" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 198475" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 198475" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 198476" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 198533" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 198533" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 198533" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 198533" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 198534" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 199289" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 199289" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 199289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 199289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 199290" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 199290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 199311" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 199311" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 199311" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 199311" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 199312" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 199379" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 199379" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 199379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 199379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 199380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 199385" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 199385" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 199385" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 199385" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 199386" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 199443" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 199443" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 199443" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 199443" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 199444" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 200199" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 200199" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 200199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 200199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 200200" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 200200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 200221" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 200221" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 200221" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 200221" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 200222" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 200289" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 200289" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 200289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 200289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 200290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 200295" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 200295" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 200295" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 200295" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 200296" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 200353" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 200353" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 200353" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 200353" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 200354" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 201109" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 201109" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 201109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 201109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 201110" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 201110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 201131" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 201131" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 201131" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 201131" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 201132" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 201199" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 201199" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 201199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 201199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 201200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 201205" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 201205" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 201205" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 201205" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 201206" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 201263" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 201263" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 201263" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 201263" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 201264" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 202019" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 202019" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 202019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 202019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 202020" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 202020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 202041" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 202041" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 202041" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 202041" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 202042" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 202109" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 202109" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 202109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 202109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 202110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 202115" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 202115" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 202115" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 202115" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 202116" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 202173" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 202173" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 202173" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 202173" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 202174" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 202929" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 202929" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 202929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 202929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 202930" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 202930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 202951" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 202951" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 202951" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 202951" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 202952" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 203019" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 203019" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 203019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 203019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 203020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 203025" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 203025" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 203025" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 203025" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 203026" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 203083" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 203083" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 203083" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 203083" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 203084" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 203839" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 203839" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 203839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 203839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 203840" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 203840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 203861" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 203861" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 203861" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 203861" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 203862" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 203929" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 203929" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 203929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 203929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 203930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 203935" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 203935" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 203935" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 203935" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 203936" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 203993" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 203993" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 203993" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 203993" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 203994" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 204749" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 204749" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 204749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 204749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 204750" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 204750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 204771" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 204771" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 204771" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 204771" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 204772" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 204839" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 204839" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 204839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 204839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 204840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 204845" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 204845" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 204845" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 204845" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 204846" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 204903" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 204903" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 204903" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 204903" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 204904" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 205659" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 205659" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 205659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 205659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 205660" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 205660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 205681" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 205681" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 205681" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 205681" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 205682" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 205749" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 205749" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 205749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 205749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 205750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 205755" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 205755" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 205755" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 205755" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 205756" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 205813" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 205813" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 205813" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 205813" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 205814" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 206569" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 206569" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 206569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 206569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 206570" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 206570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 206591" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 206591" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 206591" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 206591" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 206592" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 206659" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 206659" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 206659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 206659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 206660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 206665" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 206665" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 206665" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 206665" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 206666" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 206723" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 206723" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 206723" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 206723" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 206724" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 207479" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 207479" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 207479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 207479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 207480" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 207480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 207501" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 207501" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 207501" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 207501" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 207502" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 207569" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 207569" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 207569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 207569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 207570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 207575" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 207575" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 207575" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 207575" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 207576" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 207633" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 207633" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 207633" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 207633" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 207634" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 208389" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 208389" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 208389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 208389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 208390" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 208390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 208411" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 208411" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 208411" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 208411" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 208412" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 208479" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 208479" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 208479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 208479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 208480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 208485" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 208485" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 208485" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 208485" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 208486" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 208543" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 208543" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 208543" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 208543" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 208544" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 209299" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 209299" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 209299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 209299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 209300" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 209300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 209321" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 209321" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 209321" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 209321" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 209322" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 209389" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 209389" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 209389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 209389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 209390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 209395" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 209395" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 209395" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 209395" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 209396" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 209453" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 209453" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 209453" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 209453" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 209454" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 210209" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 210209" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 210209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 210209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 210210" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 210210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 210231" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 210231" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 210231" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 210231" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 210232" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 210299" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 210299" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 210299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 210299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 210300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 210305" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 210305" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 210305" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 210305" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 210306" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 210363" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 210363" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 210363" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 210363" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 210364" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 211119" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 211119" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 211119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 211119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 211120" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 211120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 211141" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 211141" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 211141" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 211141" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 211142" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 211209" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 211209" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 211209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 211209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 211210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 211215" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 211215" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 211215" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 211215" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 211216" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 211273" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 211273" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 211273" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 211273" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 211274" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 212029" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 212029" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 212029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 212029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 212030" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 212030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 212051" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 212051" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 212051" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 212051" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 212052" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 212119" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 212119" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 212119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 212119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 212120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 212125" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 212125" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 212125" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 212125" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 212126" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 212183" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 212183" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 212183" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 212183" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 212184" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 212939" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 212939" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 212939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 212939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 212940" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 212940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 212961" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 212961" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 212961" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 212961" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 212962" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 213029" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 213029" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 213029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 213029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 213030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 213035" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 213035" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 213035" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 213035" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 213036" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 213093" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 213093" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 213093" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 213093" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 213094" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 213849" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 213849" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 213849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 213849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 213850" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 213850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 213871" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 213871" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 213871" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 213871" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 213872" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 213939" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 213939" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 213939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 213939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 213940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 213945" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 213945" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 213945" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 213945" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 213946" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 214003" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 214003" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 214003" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 214003" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 214004" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 214759" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 214759" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 214759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 214759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 214760" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 214760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 214781" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 214781" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 214781" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 214781" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 214782" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 214849" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 214849" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 214849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 214849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 214850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 214855" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 214855" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 214855" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 214855" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 214856" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 214913" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 214913" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 214913" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 214913" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 214914" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 215669" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 215669" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 215669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 215669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 215670" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 215670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 215691" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 215691" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 215691" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 215691" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 215692" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 215759" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 215759" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 215759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 215759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 215760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 215765" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 215765" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 215765" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 215765" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 215766" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 215823" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 215823" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 215823" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 215823" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 215824" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 216579" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 216579" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 216579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 216579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 216580" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 216580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 216601" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 216601" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 216601" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 216601" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 216602" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 216669" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 216669" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 216669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 216669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 216670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 216675" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 216675" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 216675" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 216675" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 216676" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 216733" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 216733" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 216733" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 216733" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 216734" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 217489" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 217489" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 217489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 217489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 217490" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 217490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 217511" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 217511" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 217511" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 217511" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 217512" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 217579" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 217579" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 217579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 217579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 217580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 217585" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 217585" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 217585" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 217585" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 217586" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 217643" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 217643" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 217643" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 217643" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 217644" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 218399" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 218399" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 218399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 218399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 218400" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 218400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 218421" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 218421" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 218421" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 218421" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 218422" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 218489" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 218489" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 218489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 218489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 218490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 218495" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 218495" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 218495" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 218495" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 218496" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 218553" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 218553" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 218553" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 218553" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 218554" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 219309" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 219309" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 219309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 219309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 219310" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 219310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 219331" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 219331" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 219331" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 219331" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 219332" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 219399" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 219399" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 219399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 219399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 219400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 219405" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 219405" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 219405" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 219405" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 219406" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 219463" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 219463" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 219463" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 219463" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 219464" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 220219" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 220219" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 220219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 220219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 220220" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 220220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 220241" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 220241" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 220241" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 220241" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 220242" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 220309" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 220309" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 220309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 220309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 220310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 220315" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 220315" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 220315" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 220315" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 220316" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 220373" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 220373" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 220373" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 220373" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 220374" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 221129" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 221129" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 221129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 221129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 221130" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 221130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 221151" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 221151" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 221151" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 221151" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 221152" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 221219" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 221219" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 221219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 221219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 221220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 221225" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 221225" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 221225" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 221225" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 221226" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 221283" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 221283" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 221283" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 221283" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 221284" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 222039" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 222039" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 222039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 222039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 222040" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 222040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 222061" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 222061" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 222061" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 222061" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 222062" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 222129" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 222129" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 222129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 222129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 222130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 222135" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 222135" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 222135" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 222135" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 222136" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 222193" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 222193" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 222193" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 222193" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 222194" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 222949" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 222949" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 222949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 222949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 222950" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 222950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 222971" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 222971" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 222971" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 222971" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 222972" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 223039" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 223039" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 223039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 223039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 223040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 223045" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 223045" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 223045" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 223045" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 223046" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 223103" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 223103" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 223103" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 223103" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 223104" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 223859" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 223859" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 223859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 223859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 223860" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 223860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 223881" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 223881" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 223881" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 223881" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 223882" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 223949" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 223949" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 223949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 223949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 223950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 223955" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 223955" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 223955" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 223955" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 223956" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 224013" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 224013" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 224013" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 224013" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 224014" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 224769" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 224769" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 224769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 224769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 224770" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 224770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 224791" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 224791" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 224791" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 224791" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 224792" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 224859" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 224859" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 224859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 224859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 224860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 224865" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 224865" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 224865" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 224865" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 224866" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 224923" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 224923" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 224923" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 224923" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 224924" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 225679" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 225679" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 225679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 225679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 225680" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 225680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 225701" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 225701" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 225701" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 225701" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 225702" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 225769" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 225769" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 225769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 225769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 225770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 225775" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 225775" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 225775" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 225775" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 225776" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 225833" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 225833" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 225833" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 225833" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 225834" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 226589" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 226589" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 226589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 226589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 226590" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 226590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 226611" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 226611" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 226611" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 226611" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 226612" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 226679" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 226679" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 226679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 226679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 226680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 226685" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 226685" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 226685" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 226685" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 226686" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 226743" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 226743" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 226743" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 226743" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 226744" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 227499" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 227499" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 227499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 227499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 227500" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 227500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 227521" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 227521" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 227521" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 227521" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 227522" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 227589" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 227589" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 227589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 227589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 227590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 227595" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 227595" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 227595" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 227595" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 227596" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 227653" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 227653" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 227653" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 227653" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 227654" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 228409" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 228409" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 228409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 228409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 228410" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 228410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 228431" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 228431" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 228431" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 228431" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 228432" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 228499" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 228499" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 228499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 228499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 228500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 228505" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 228505" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 228505" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 228505" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 228506" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 228563" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 228563" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 228563" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 228563" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 228564" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 229319" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 229319" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 229319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 229319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 229320" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 229320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 229341" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 229341" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 229341" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 229341" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 229342" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 229409" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 229409" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 229409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 229409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 229410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 229415" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 229415" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 229415" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 229415" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 229416" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 229473" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 229473" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 229473" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 229473" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 229474" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 230229" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 230229" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 230229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 230229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 230230" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 230230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 230251" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 230251" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 230251" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 230251" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 230252" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 230319" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 230319" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 230319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 230319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 230320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 230325" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 230325" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 230325" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 230325" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 230326" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 230383" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 230383" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 230383" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 230383" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 230384" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 231139" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 231139" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 231139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 231139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 231140" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 231140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 231161" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 231161" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 231161" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 231161" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 231162" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 231229" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 231229" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 231229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 231229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 231230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 231235" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 231235" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 231235" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 231235" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 231236" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 231293" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 231293" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 231293" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 231293" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 231294" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 232049" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 232049" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 232049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 232049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 232050" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 232050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 232071" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 232071" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 232071" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 232071" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 232072" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 232139" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 232139" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 232139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 232139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 232140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 232145" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 232145" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 232145" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 232145" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 232146" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 232203" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 232203" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 232203" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 232203" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 232204" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 232959" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 232959" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 232959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 232959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 232960" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 232960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 232981" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 232981" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 232981" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 232981" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 232982" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 233049" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 233049" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 233049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 233049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 233050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 233055" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 233055" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 233055" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 233055" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 233056" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 233113" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 233113" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 233113" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 233113" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 233114" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 233869" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 233869" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 233869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 233869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 233870" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 233870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 233891" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 233891" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 233891" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 233891" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 233892" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 233959" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 233959" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 233959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 233959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 233960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 233965" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 233965" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 233965" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 233965" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 233966" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 234023" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 234023" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 234023" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 234023" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 234024" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 234779" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 234779" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 234779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 234779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 234780" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 234780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 234801" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 234801" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 234801" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 234801" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 234802" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 234869" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 234869" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 234869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 234869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 234870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 234875" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 234875" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 234875" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 234875" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 234876" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 234933" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 234933" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 234933" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 234933" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 234934" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 235689" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 235689" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 235689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 235689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 235690" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 235690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 235711" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 235711" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 235711" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 235711" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 235712" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 235779" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 235779" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 235779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 235779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 235780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 235785" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 235785" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 235785" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 235785" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 235786" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 235843" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 235843" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 235843" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 235843" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 235844" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 236599" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 236599" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 236599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 236599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 236600" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 236600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 236621" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 236621" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 236621" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 236621" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 236622" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 236689" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 236689" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 236689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 236689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 236690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 236695" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 236695" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 236695" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 236695" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 236696" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 236753" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 236753" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 236753" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 236753" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 236754" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 237509" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 237509" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 237509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 237509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 237510" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 237510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 237531" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 237531" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 237531" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 237531" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 237532" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 237599" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 237599" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 237599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 237599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 237600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 237605" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 237605" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 237605" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 237605" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 237606" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 237663" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 237663" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 237663" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 237663" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 237664" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 238419" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 238419" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 238419" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 238419" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 238420" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 238420" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 238441" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 238441" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 238441" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 238441" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 238442" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 238509" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 238509" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 238509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 238509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 238510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 238515" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 238515" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 238515" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 238515" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 238516" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 238573" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 238573" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 238573" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 238573" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 238574" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 300);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 238874" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 238874" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 238874" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 238874" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 238875" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 238875" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 238896" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 238896" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 238896" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 238896" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 238897" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 238928" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 238928" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 238928" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 238928" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 238929" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 239329" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 239329" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 239329" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 239329" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 239330" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 239351" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 239351" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 239351" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 239351" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 239352" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 239383" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 239383" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 239383" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 239383" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 239384" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 239425" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 239425" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 239425" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 239425" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 239426" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 239806" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 239806" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 239806" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 239806" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 239807" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 239838" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 239838" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 239838" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 239838" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 239839" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 240239" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 240239" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 240239" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 240239" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 240240" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 240261" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 240261" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 240261" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 240261" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 240262" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 240293" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 240293" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 240293" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 240293" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 240294" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 240335" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 240335" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 240335" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 240335" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 240336" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 240716" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 240716" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 240716" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 240716" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 240717" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 240748" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 240748" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 240748" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 240748" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 240749" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 241149" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 241149" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 241149" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 241149" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 241150" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 241171" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 241171" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 241171" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 241171" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 241172" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 241203" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 241203" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 241203" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 241203" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 241204" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 241245" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 241245" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 241245" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 241245" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 241246" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 241626" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 241626" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 241626" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 241626" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 241627" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 386);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 242013" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 242013" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 242013" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 242013" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 242014" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 45);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 242059" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 242059" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 242059" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 242059" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 242060" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 242081" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 242081" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 242081" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 242081" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 242082" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 73);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 242155" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 242155" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 242155" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 242155" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 242156" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 312);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 242468" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 242468" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 242468" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 242468" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 242469" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 242536" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 242536" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 242536" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 242536" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 242537" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 386);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 242923" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 242923" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 242923" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 242923" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 242924" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 45);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 242969" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 242969" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 242969" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 242969" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 242970" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 242991" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 242991" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 242991" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 242991" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 242992" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 73);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 243065" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 243065" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 243065" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 243065" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 243066" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 312);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 243378" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 243378" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 243378" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 243378" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 243379" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 243446" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 243446" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 243446" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 243446" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 243447" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 386);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 243833" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 243833" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 243833" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 243833" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 243834" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 45);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 243879" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 243879" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 243879" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 243879" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 243880" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 243901" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 243901" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 243901" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 243901" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 243902" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 73);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 243975" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 243975" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 243975" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 243975" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 243976" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 312);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 244288" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 244288" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 244288" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 244288" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 244289" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 244356" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 244356" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 244356" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 244356" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 244357" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 244388" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 244388" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 244388" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 244388" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 244389" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 244789" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 244789" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 244789" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 244789" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 244790" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 244811" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 244811" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 244811" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 244811" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 244812" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 244843" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 244843" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 244843" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 244843" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 244844" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 244885" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 244885" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 244885" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 244885" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 244886" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 245266" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 245266" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 245266" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 245266" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 245267" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 245298" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 245298" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 245298" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 245298" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 245299" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 245699" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 245699" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 245699" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 245699" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 245700" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 245721" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 245721" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 245721" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 245721" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 245722" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 245753" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 245753" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 245753" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 245753" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 245754" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 245795" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 245795" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 245795" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 245795" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 245796" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 380);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 246176" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 246176" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 246176" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 246176" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 246177" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 246208" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 246208" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 246208" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 246208" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 246209" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 400);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 246609" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 246609" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 246609" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 246609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 246610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 246631" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 246631" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 246631" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 246631" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 246632" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 31);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 246663" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 246663" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 246663" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 246663" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 246664" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 41);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 246705" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 246705" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 246705" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 246705" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 246706" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 358);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 247064" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 247064" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 247064" severity error;
		assert (vsync2_prime = '0') report "Unexpected value for vsync2_prime at cycle 247064" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 247065" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 454);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 247519" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 247519" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 247519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 247519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 247520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 247541" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 247541" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 247541" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 247541" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 247542" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 247609" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 247609" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 247609" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 247609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 247610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 247615" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 247615" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 247615" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 247615" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 247616" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 248429" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 248429" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 248429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 248429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 248430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 248451" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 248451" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 248451" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 248451" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 248452" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 248519" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 248519" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 248519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 248519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 248520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 248525" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 248525" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 248525" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 248525" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 248526" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 249339" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 249339" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 249339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 249339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 249340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 249361" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 249361" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 249361" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 249361" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 249362" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 249429" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 249429" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 249429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 249429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 249430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 249435" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 249435" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 249435" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 249435" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 249436" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 250249" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 250249" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 250249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 250249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 250250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 250271" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 250271" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 250271" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 250271" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 250272" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 250339" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 250339" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 250339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 250339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 250340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 250345" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 250345" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 250345" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 250345" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 250346" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 251159" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 251159" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 251159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 251159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 251160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 251181" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 251181" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 251181" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 251181" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 251182" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 251249" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 251249" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 251249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 251249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 251250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 251255" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 251255" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 251255" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 251255" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 251256" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 252069" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 252069" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 252069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 252069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 252070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 252091" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 252091" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 252091" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 252091" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 252092" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 252159" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 252159" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 252159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 252159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 252160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 252165" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 252165" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 252165" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 252165" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 252166" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 252979" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 252979" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 252979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 252979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 252980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 253001" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 253001" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 253001" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 253001" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 253002" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 253069" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 253069" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 253069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 253069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 253070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 253075" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 253075" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 253075" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 253075" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 253076" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 253889" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 253889" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 253889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 253889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 253890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 253911" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 253911" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 253911" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 253911" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 253912" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 253979" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 253979" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 253979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 253979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 253980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 253985" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 253985" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 253985" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 253985" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 253986" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 254799" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 254799" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 254799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 254799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 254800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 254821" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 254821" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 254821" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 254821" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 254822" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 254889" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 254889" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 254889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 254889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 254890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 254895" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 254895" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 254895" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 254895" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 254896" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 255709" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 255709" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 255709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 255709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 255710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 255731" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 255731" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 255731" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 255731" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 255732" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 255799" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 255799" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 255799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 255799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 255800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 255805" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 255805" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 255805" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 255805" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 255806" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 813);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 256619" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 256619" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 256619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 256619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 256620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 256641" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 256641" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 256641" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 256641" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 256642" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 256709" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 256709" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 256709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 256709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 256710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 256715" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 256715" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 256715" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 256715" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 256716" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 512);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 257228" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 257228" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 257228" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 257228" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 257229" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 300);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 257529" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 257529" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 257529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 257529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 257530" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 257530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 257551" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 257551" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 257551" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 257551" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 257552" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 257619" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 257619" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 257619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 257619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 257620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 257625" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 257625" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 257625" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 257625" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 257626" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 257683" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 257683" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 257683" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 257683" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 257684" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 258439" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 258439" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 258439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 258439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 258440" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 258440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 258461" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 258461" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 258461" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 258461" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 258462" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 258529" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 258529" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 258529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 258529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 258530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 258535" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 258535" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 258535" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 258535" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 258536" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 258593" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 258593" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 258593" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 258593" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 258594" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 259349" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 259349" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 259349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 259349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 259350" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 259350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 259371" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 259371" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 259371" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 259371" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 259372" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 259439" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 259439" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 259439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 259439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 259440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 259445" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 259445" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 259445" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 259445" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 259446" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 259503" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 259503" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 259503" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 259503" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 259504" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 260259" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 260259" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 260259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 260259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 260260" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 260260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 260281" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 260281" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 260281" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 260281" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 260282" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 260349" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 260349" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 260349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 260349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 260350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 260355" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 260355" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 260355" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 260355" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 260356" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 260413" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 260413" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 260413" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 260413" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 260414" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 261169" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 261169" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 261169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 261169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 261170" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 261170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 261191" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 261191" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 261191" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 261191" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 261192" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 261259" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 261259" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 261259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 261259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 261260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 261265" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 261265" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 261265" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 261265" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 261266" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 261323" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 261323" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 261323" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 261323" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 261324" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 262079" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 262079" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 262079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 262079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 262080" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 262080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 262101" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 262101" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 262101" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 262101" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 262102" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 262169" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 262169" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 262169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 262169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 262170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 262175" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 262175" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 262175" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 262175" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 262176" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 262233" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 262233" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 262233" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 262233" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 262234" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 262989" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 262989" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 262989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 262989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 262990" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 262990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 263011" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 263011" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 263011" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 263011" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 263012" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 263079" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 263079" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 263079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 263079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 263080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 263085" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 263085" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 263085" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 263085" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 263086" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 263143" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 263143" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 263143" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 263143" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 263144" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 263899" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 263899" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 263899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 263899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 263900" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 263900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 263921" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 263921" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 263921" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 263921" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 263922" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 263989" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 263989" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 263989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 263989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 263990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 263995" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 263995" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 263995" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 263995" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 263996" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 264053" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 264053" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 264053" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 264053" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 264054" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 264809" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 264809" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 264809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 264809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 264810" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 264810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 264831" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 264831" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 264831" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 264831" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 264832" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 264899" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 264899" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 264899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 264899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 264900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 264905" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 264905" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 264905" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 264905" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 264906" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 264963" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 264963" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 264963" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 264963" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 264964" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 265719" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 265719" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 265719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 265719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 265720" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 265720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 265741" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 265741" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 265741" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 265741" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 265742" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 265809" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 265809" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 265809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 265809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 265810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 265815" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 265815" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 265815" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 265815" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 265816" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 265873" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 265873" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 265873" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 265873" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 265874" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 266629" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 266629" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 266629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 266629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 266630" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 266630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 266651" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 266651" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 266651" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 266651" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 266652" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 266719" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 266719" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 266719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 266719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 266720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 266725" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 266725" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 266725" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 266725" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 266726" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 266783" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 266783" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 266783" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 266783" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 266784" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 267539" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 267539" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 267539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 267539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 267540" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 267540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 267561" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 267561" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 267561" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 267561" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 267562" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 267629" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 267629" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 267629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 267629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 267630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 267635" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 267635" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 267635" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 267635" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 267636" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 267693" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 267693" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 267693" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 267693" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 267694" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 268449" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 268449" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 268449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 268449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 268450" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 268450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 268471" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 268471" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 268471" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 268471" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 268472" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 268539" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 268539" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 268539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 268539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 268540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 268545" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 268545" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 268545" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 268545" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 268546" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 268603" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 268603" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 268603" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 268603" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 268604" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 269359" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 269359" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 269359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 269359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 269360" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 269360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 269381" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 269381" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 269381" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 269381" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 269382" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 269449" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 269449" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 269449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 269449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 269450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 269455" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 269455" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 269455" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 269455" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 269456" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 269513" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 269513" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 269513" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 269513" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 269514" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 270269" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 270269" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 270269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 270269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 270270" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 270270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 270291" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 270291" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 270291" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 270291" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 270292" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 270359" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 270359" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 270359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 270359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 270360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 270365" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 270365" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 270365" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 270365" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 270366" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 270423" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 270423" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 270423" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 270423" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 270424" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 271179" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 271179" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 271179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 271179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 271180" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 271180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 271201" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 271201" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 271201" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 271201" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 271202" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 271269" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 271269" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 271269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 271269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 271270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 271275" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 271275" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 271275" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 271275" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 271276" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 271333" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 271333" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 271333" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 271333" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 271334" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 272089" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 272089" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 272089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 272089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 272090" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 272090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 272111" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 272111" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 272111" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 272111" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 272112" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 272179" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 272179" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 272179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 272179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 272180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 272185" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 272185" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 272185" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 272185" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 272186" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 272243" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 272243" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 272243" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 272243" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 272244" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 272999" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 272999" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 272999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 272999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 273000" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 273000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 273021" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 273021" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 273021" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 273021" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 273022" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 273089" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 273089" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 273089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 273089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 273090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 273095" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 273095" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 273095" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 273095" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 273096" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 273153" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 273153" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 273153" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 273153" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 273154" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 273909" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 273909" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 273909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 273909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 273910" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 273910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 273931" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 273931" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 273931" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 273931" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 273932" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 273999" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 273999" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 273999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 273999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 274000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 274005" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 274005" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 274005" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 274005" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 274006" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 274063" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 274063" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 274063" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 274063" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 274064" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 274819" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 274819" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 274819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 274819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 274820" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 274820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 274841" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 274841" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 274841" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 274841" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 274842" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 274909" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 274909" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 274909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 274909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 274910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 274915" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 274915" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 274915" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 274915" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 274916" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 274973" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 274973" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 274973" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 274973" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 274974" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 275729" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 275729" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 275729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 275729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 275730" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 275730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 275751" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 275751" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 275751" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 275751" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 275752" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 275819" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 275819" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 275819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 275819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 275820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 275825" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 275825" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 275825" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 275825" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 275826" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 275883" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 275883" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 275883" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 275883" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 275884" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 276639" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 276639" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 276639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 276639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 276640" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 276640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 276661" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 276661" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 276661" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 276661" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 276662" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 276729" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 276729" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 276729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 276729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 276730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 276735" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 276735" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 276735" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 276735" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 276736" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 276793" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 276793" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 276793" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 276793" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 276794" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 277549" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 277549" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 277549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 277549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 277550" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 277550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 277571" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 277571" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 277571" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 277571" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 277572" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 277639" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 277639" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 277639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 277639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 277640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 277645" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 277645" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 277645" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 277645" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 277646" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 277703" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 277703" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 277703" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 277703" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 277704" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 278459" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 278459" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 278459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 278459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 278460" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 278460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 278481" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 278481" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 278481" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 278481" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 278482" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 278549" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 278549" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 278549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 278549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 278550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 278555" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 278555" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 278555" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 278555" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 278556" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 278613" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 278613" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 278613" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 278613" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 278614" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 279369" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 279369" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 279369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 279369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 279370" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 279370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 279391" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 279391" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 279391" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 279391" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 279392" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 279459" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 279459" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 279459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 279459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 279460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 279465" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 279465" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 279465" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 279465" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 279466" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 279523" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 279523" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 279523" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 279523" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 279524" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 280279" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 280279" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 280279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 280279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 280280" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 280280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 280301" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 280301" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 280301" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 280301" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 280302" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 280369" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 280369" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 280369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 280369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 280370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 280375" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 280375" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 280375" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 280375" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 280376" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 280433" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 280433" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 280433" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 280433" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 280434" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 281189" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 281189" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 281189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 281189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 281190" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 281190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 281211" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 281211" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 281211" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 281211" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 281212" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 281279" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 281279" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 281279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 281279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 281280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 281285" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 281285" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 281285" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 281285" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 281286" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 281343" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 281343" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 281343" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 281343" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 281344" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 282099" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 282099" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 282099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 282099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 282100" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 282100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 282121" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 282121" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 282121" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 282121" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 282122" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 282189" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 282189" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 282189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 282189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 282190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 282195" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 282195" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 282195" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 282195" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 282196" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 282253" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 282253" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 282253" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 282253" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 282254" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 283009" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 283009" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 283009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 283009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 283010" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 283010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 283031" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 283031" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 283031" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 283031" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 283032" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 283099" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 283099" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 283099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 283099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 283100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 283105" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 283105" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 283105" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 283105" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 283106" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 283163" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 283163" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 283163" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 283163" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 283164" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 283919" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 283919" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 283919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 283919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 283920" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 283920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 283941" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 283941" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 283941" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 283941" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 283942" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 284009" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 284009" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 284009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 284009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 284010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 284015" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 284015" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 284015" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 284015" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 284016" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 284073" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 284073" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 284073" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 284073" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 284074" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 284829" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 284829" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 284829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 284829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 284830" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 284830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 284851" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 284851" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 284851" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 284851" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 284852" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 284919" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 284919" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 284919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 284919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 284920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 284925" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 284925" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 284925" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 284925" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 284926" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 284983" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 284983" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 284983" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 284983" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 284984" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 285739" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 285739" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 285739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 285739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 285740" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 285740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 285761" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 285761" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 285761" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 285761" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 285762" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 285829" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 285829" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 285829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 285829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 285830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 285835" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 285835" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 285835" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 285835" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 285836" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 285893" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 285893" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 285893" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 285893" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 285894" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 286649" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 286649" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 286649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 286649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 286650" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 286650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 286671" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 286671" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 286671" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 286671" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 286672" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 286739" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 286739" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 286739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 286739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 286740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 286745" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 286745" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 286745" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 286745" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 286746" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 286803" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 286803" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 286803" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 286803" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 286804" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 287559" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 287559" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 287559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 287559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 287560" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 287560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 287581" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 287581" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 287581" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 287581" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 287582" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 287649" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 287649" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 287649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 287649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 287650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 287655" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 287655" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 287655" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 287655" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 287656" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 287713" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 287713" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 287713" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 287713" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 287714" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 288469" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 288469" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 288469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 288469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 288470" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 288470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 288491" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 288491" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 288491" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 288491" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 288492" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 288559" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 288559" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 288559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 288559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 288560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 288565" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 288565" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 288565" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 288565" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 288566" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 288623" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 288623" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 288623" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 288623" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 288624" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 289379" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 289379" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 289379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 289379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 289380" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 289380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 289401" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 289401" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 289401" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 289401" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 289402" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 289469" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 289469" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 289469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 289469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 289470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 289475" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 289475" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 289475" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 289475" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 289476" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 289533" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 289533" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 289533" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 289533" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 289534" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 290289" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 290289" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 290289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 290289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 290290" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 290290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 290311" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 290311" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 290311" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 290311" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 290312" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 290379" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 290379" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 290379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 290379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 290380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 290385" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 290385" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 290385" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 290385" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 290386" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 290443" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 290443" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 290443" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 290443" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 290444" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 291199" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 291199" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 291199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 291199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 291200" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 291200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 291221" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 291221" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 291221" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 291221" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 291222" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 291289" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 291289" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 291289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 291289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 291290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 291295" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 291295" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 291295" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 291295" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 291296" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 291353" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 291353" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 291353" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 291353" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 291354" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 292109" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 292109" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 292109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 292109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 292110" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 292110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 292131" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 292131" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 292131" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 292131" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 292132" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 292199" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 292199" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 292199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 292199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 292200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 292205" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 292205" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 292205" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 292205" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 292206" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 292263" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 292263" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 292263" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 292263" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 292264" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 293019" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 293019" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 293019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 293019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 293020" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 293020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 293041" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 293041" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 293041" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 293041" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 293042" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 293109" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 293109" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 293109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 293109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 293110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 293115" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 293115" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 293115" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 293115" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 293116" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 293173" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 293173" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 293173" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 293173" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 293174" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 293929" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 293929" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 293929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 293929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 293930" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 293930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 293951" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 293951" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 293951" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 293951" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 293952" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 294019" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 294019" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 294019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 294019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 294020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 294025" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 294025" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 294025" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 294025" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 294026" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 294083" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 294083" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 294083" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 294083" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 294084" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 294839" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 294839" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 294839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 294839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 294840" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 294840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 294861" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 294861" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 294861" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 294861" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 294862" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 294929" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 294929" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 294929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 294929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 294930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 294935" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 294935" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 294935" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 294935" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 294936" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 294993" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 294993" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 294993" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 294993" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 294994" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 295749" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 295749" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 295749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 295749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 295750" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 295750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 295771" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 295771" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 295771" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 295771" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 295772" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 295839" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 295839" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 295839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 295839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 295840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 295845" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 295845" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 295845" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 295845" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 295846" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 295903" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 295903" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 295903" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 295903" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 295904" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 296659" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 296659" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 296659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 296659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 296660" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 296660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 296681" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 296681" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 296681" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 296681" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 296682" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 296749" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 296749" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 296749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 296749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 296750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 296755" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 296755" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 296755" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 296755" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 296756" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 296813" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 296813" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 296813" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 296813" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 296814" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 297569" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 297569" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 297569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 297569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 297570" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 297570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 297591" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 297591" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 297591" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 297591" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 297592" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 297659" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 297659" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 297659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 297659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 297660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 297665" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 297665" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 297665" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 297665" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 297666" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 297723" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 297723" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 297723" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 297723" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 297724" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 298479" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 298479" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 298479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 298479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 298480" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 298480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 298501" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 298501" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 298501" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 298501" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 298502" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 298569" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 298569" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 298569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 298569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 298570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 298575" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 298575" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 298575" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 298575" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 298576" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 298633" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 298633" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 298633" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 298633" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 298634" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 299389" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 299389" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 299389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 299389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 299390" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 299390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 299411" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 299411" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 299411" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 299411" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 299412" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 299479" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 299479" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 299479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 299479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 299480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 299485" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 299485" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 299485" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 299485" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 299486" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 299543" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 299543" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 299543" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 299543" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 299544" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 300299" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 300299" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 300299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 300299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 300300" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 300300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 300321" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 300321" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 300321" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 300321" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 300322" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 300389" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 300389" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 300389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 300389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 300390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 300395" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 300395" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 300395" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 300395" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 300396" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 300453" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 300453" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 300453" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 300453" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 300454" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 301209" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 301209" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 301209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 301209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 301210" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 301210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 301231" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 301231" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 301231" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 301231" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 301232" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 301299" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 301299" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 301299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 301299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 301300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 301305" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 301305" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 301305" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 301305" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 301306" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 301363" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 301363" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 301363" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 301363" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 301364" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 302119" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 302119" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 302119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 302119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 302120" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 302120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 302141" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 302141" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 302141" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 302141" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 302142" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 302209" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 302209" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 302209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 302209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 302210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 302215" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 302215" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 302215" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 302215" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 302216" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 302273" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 302273" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 302273" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 302273" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 302274" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 303029" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 303029" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 303029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 303029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 303030" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 303030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 303051" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 303051" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 303051" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 303051" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 303052" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 303119" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 303119" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 303119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 303119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 303120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 303125" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 303125" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 303125" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 303125" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 303126" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 303183" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 303183" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 303183" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 303183" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 303184" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 303939" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 303939" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 303939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 303939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 303940" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 303940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 303961" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 303961" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 303961" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 303961" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 303962" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 304029" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 304029" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 304029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 304029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 304030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 304035" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 304035" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 304035" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 304035" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 304036" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 304093" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 304093" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 304093" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 304093" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 304094" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 304849" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 304849" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 304849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 304849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 304850" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 304850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 304871" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 304871" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 304871" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 304871" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 304872" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 304939" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 304939" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 304939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 304939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 304940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 304945" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 304945" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 304945" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 304945" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 304946" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 305003" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 305003" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 305003" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 305003" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 305004" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 305759" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 305759" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 305759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 305759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 305760" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 305760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 305781" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 305781" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 305781" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 305781" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 305782" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 305849" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 305849" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 305849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 305849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 305850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 305855" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 305855" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 305855" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 305855" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 305856" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 305913" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 305913" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 305913" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 305913" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 305914" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 306669" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 306669" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 306669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 306669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 306670" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 306670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 306691" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 306691" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 306691" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 306691" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 306692" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 306759" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 306759" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 306759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 306759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 306760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 306765" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 306765" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 306765" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 306765" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 306766" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 306823" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 306823" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 306823" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 306823" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 306824" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 307579" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 307579" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 307579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 307579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 307580" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 307580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 307601" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 307601" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 307601" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 307601" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 307602" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 307669" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 307669" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 307669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 307669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 307670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 307675" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 307675" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 307675" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 307675" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 307676" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 307733" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 307733" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 307733" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 307733" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 307734" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 308489" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 308489" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 308489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 308489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 308490" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 308490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 308511" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 308511" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 308511" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 308511" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 308512" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 308579" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 308579" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 308579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 308579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 308580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 308585" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 308585" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 308585" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 308585" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 308586" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 308643" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 308643" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 308643" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 308643" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 308644" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 309399" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 309399" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 309399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 309399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 309400" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 309400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 309421" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 309421" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 309421" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 309421" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 309422" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 309489" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 309489" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 309489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 309489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 309490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 309495" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 309495" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 309495" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 309495" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 309496" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 309553" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 309553" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 309553" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 309553" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 309554" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 310309" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 310309" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 310309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 310309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 310310" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 310310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 310331" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 310331" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 310331" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 310331" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 310332" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 310399" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 310399" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 310399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 310399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 310400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 310405" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 310405" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 310405" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 310405" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 310406" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 310463" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 310463" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 310463" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 310463" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 310464" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 311219" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 311219" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 311219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 311219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 311220" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 311220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 311241" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 311241" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 311241" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 311241" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 311242" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 311309" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 311309" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 311309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 311309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 311310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 311315" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 311315" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 311315" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 311315" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 311316" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 311373" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 311373" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 311373" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 311373" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 311374" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 312129" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 312129" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 312129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 312129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 312130" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 312130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 312151" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 312151" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 312151" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 312151" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 312152" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 312219" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 312219" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 312219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 312219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 312220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 312225" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 312225" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 312225" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 312225" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 312226" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 312283" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 312283" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 312283" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 312283" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 312284" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 313039" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 313039" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 313039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 313039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 313040" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 313040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 313061" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 313061" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 313061" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 313061" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 313062" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 313129" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 313129" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 313129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 313129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 313130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 313135" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 313135" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 313135" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 313135" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 313136" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 313193" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 313193" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 313193" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 313193" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 313194" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 313949" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 313949" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 313949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 313949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 313950" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 313950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 313971" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 313971" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 313971" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 313971" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 313972" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 314039" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 314039" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 314039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 314039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 314040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 314045" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 314045" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 314045" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 314045" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 314046" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 314103" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 314103" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 314103" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 314103" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 314104" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 314859" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 314859" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 314859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 314859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 314860" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 314860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 314881" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 314881" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 314881" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 314881" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 314882" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 314949" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 314949" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 314949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 314949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 314950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 314955" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 314955" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 314955" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 314955" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 314956" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 315013" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 315013" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 315013" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 315013" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 315014" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 315769" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 315769" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 315769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 315769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 315770" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 315770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 315791" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 315791" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 315791" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 315791" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 315792" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 315859" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 315859" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 315859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 315859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 315860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 315865" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 315865" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 315865" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 315865" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 315866" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 315923" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 315923" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 315923" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 315923" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 315924" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 316679" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 316679" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 316679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 316679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 316680" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 316680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 316701" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 316701" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 316701" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 316701" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 316702" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 316769" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 316769" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 316769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 316769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 316770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 316775" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 316775" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 316775" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 316775" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 316776" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 316833" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 316833" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 316833" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 316833" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 316834" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 317589" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 317589" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 317589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 317589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 317590" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 317590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 317611" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 317611" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 317611" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 317611" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 317612" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 317679" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 317679" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 317679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 317679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 317680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 317685" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 317685" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 317685" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 317685" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 317686" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 317743" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 317743" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 317743" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 317743" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 317744" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 318499" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 318499" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 318499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 318499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 318500" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 318500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 318521" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 318521" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 318521" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 318521" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 318522" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 318589" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 318589" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 318589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 318589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 318590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 318595" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 318595" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 318595" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 318595" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 318596" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 318653" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 318653" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 318653" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 318653" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 318654" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 319409" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 319409" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 319409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 319409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 319410" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 319410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 319431" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 319431" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 319431" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 319431" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 319432" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 319499" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 319499" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 319499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 319499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 319500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 319505" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 319505" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 319505" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 319505" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 319506" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 319563" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 319563" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 319563" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 319563" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 319564" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 320319" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 320319" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 320319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 320319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 320320" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 320320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 320341" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 320341" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 320341" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 320341" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 320342" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 320409" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 320409" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 320409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 320409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 320410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 320415" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 320415" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 320415" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 320415" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 320416" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 320473" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 320473" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 320473" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 320473" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 320474" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 321229" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 321229" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 321229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 321229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 321230" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 321230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 321251" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 321251" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 321251" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 321251" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 321252" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 321319" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 321319" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 321319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 321319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 321320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 321325" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 321325" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 321325" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 321325" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 321326" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 321383" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 321383" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 321383" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 321383" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 321384" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 322139" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 322139" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 322139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 322139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 322140" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 322140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 322161" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 322161" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 322161" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 322161" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 322162" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 322229" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 322229" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 322229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 322229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 322230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 322235" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 322235" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 322235" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 322235" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 322236" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 322293" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 322293" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 322293" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 322293" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 322294" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 323049" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 323049" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 323049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 323049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 323050" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 323050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 323071" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 323071" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 323071" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 323071" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 323072" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 323139" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 323139" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 323139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 323139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 323140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 323145" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 323145" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 323145" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 323145" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 323146" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 323203" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 323203" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 323203" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 323203" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 323204" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 323959" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 323959" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 323959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 323959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 323960" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 323960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 323981" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 323981" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 323981" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 323981" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 323982" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 324049" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 324049" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 324049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 324049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 324050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 324055" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 324055" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 324055" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 324055" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 324056" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 324113" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 324113" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 324113" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 324113" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 324114" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 324869" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 324869" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 324869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 324869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 324870" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 324870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 324891" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 324891" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 324891" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 324891" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 324892" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 324959" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 324959" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 324959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 324959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 324960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 324965" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 324965" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 324965" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 324965" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 324966" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 325023" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 325023" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 325023" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 325023" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 325024" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 325779" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 325779" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 325779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 325779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 325780" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 325780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 325801" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 325801" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 325801" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 325801" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 325802" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 325869" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 325869" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 325869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 325869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 325870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 325875" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 325875" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 325875" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 325875" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 325876" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 325933" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 325933" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 325933" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 325933" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 325934" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 326689" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 326689" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 326689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 326689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 326690" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 326690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 326711" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 326711" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 326711" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 326711" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 326712" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 326779" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 326779" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 326779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 326779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 326780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 326785" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 326785" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 326785" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 326785" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 326786" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 326843" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 326843" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 326843" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 326843" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 326844" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 327599" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 327599" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 327599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 327599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 327600" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 327600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 327621" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 327621" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 327621" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 327621" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 327622" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 327689" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 327689" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 327689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 327689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 327690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 327695" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 327695" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 327695" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 327695" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 327696" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 327753" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 327753" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 327753" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 327753" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 327754" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 328509" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 328509" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 328509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 328509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 328510" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 328510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 328531" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 328531" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 328531" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 328531" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 328532" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 328599" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 328599" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 328599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 328599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 328600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 328605" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 328605" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 328605" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 328605" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 328606" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 328663" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 328663" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 328663" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 328663" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 328664" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 329419" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 329419" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 329419" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 329419" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 329420" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 329420" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 329441" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 329441" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 329441" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 329441" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 329442" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 329509" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 329509" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 329509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 329509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 329510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 329515" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 329515" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 329515" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 329515" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 329516" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 329573" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 329573" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 329573" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 329573" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 329574" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 330329" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 330329" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 330329" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 330329" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 330330" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 330330" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 330351" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 330351" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 330351" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 330351" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 330352" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 330419" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 330419" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 330419" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 330419" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 330420" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 330425" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 330425" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 330425" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 330425" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 330426" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 330483" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 330483" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 330483" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 330483" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 330484" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 331239" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 331239" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 331239" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 331239" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 331240" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 331240" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 331261" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 331261" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 331261" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 331261" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 331262" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 331329" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 331329" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 331329" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 331329" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 331330" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 331335" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 331335" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 331335" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 331335" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 331336" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 331393" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 331393" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 331393" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 331393" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 331394" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 332149" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 332149" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 332149" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 332149" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 332150" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 332150" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 332171" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 332171" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 332171" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 332171" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 332172" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 332239" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 332239" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 332239" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 332239" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 332240" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 332245" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 332245" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 332245" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 332245" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 332246" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 332303" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 332303" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 332303" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 332303" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 332304" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 333059" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 333059" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 333059" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 333059" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 333060" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 333060" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 333081" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 333081" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 333081" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 333081" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 333082" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 333149" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 333149" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 333149" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 333149" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 333150" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 333155" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 333155" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 333155" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 333155" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 333156" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 333213" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 333213" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 333213" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 333213" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 333214" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 333969" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 333969" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 333969" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 333969" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 333970" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 333970" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 333991" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 333991" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 333991" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 333991" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 333992" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 334059" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 334059" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 334059" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 334059" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 334060" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 334065" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 334065" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 334065" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 334065" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 334066" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 334123" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 334123" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 334123" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 334123" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 334124" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 334879" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 334879" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 334879" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 334879" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 334880" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 334880" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 334901" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 334901" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 334901" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 334901" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 334902" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 334969" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 334969" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 334969" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 334969" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 334970" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 334975" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 334975" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 334975" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 334975" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 334976" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 335033" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 335033" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 335033" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 335033" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 335034" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 335789" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 335789" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 335789" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 335789" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 335790" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 335790" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 335811" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 335811" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 335811" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 335811" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 335812" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 335879" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 335879" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 335879" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 335879" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 335880" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 335885" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 335885" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 335885" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 335885" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 335886" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 335943" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 335943" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 335943" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 335943" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 335944" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 336699" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 336699" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 336699" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 336699" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 336700" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 336700" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 336721" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 336721" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 336721" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 336721" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 336722" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 336789" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 336789" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 336789" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 336789" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 336790" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 336795" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 336795" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 336795" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 336795" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 336796" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 336853" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 336853" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 336853" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 336853" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 336854" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 337609" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 337609" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 337609" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 337609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 337610" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 337610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 337631" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 337631" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 337631" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 337631" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 337632" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 337699" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 337699" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 337699" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 337699" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 337700" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 337705" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 337705" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 337705" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 337705" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 337706" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 337763" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 337763" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 337763" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 337763" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 337764" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 338519" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 338519" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 338519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 338519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 338520" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 338520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 338541" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 338541" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 338541" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 338541" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 338542" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 338609" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 338609" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 338609" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 338609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 338610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 338615" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 338615" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 338615" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 338615" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 338616" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 338673" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 338673" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 338673" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 338673" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 338674" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 339429" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 339429" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 339429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 339429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 339430" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 339430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 339451" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 339451" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 339451" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 339451" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 339452" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 339519" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 339519" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 339519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 339519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 339520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 339525" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 339525" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 339525" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 339525" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 339526" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 339583" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 339583" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 339583" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 339583" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 339584" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 340339" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 340339" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 340339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 340339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 340340" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 340340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 340361" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 340361" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 340361" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 340361" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 340362" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 340429" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 340429" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 340429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 340429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 340430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 340435" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 340435" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 340435" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 340435" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 340436" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 340493" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 340493" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 340493" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 340493" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 340494" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 341249" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 341249" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 341249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 341249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 341250" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 341250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 341271" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 341271" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 341271" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 341271" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 341272" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 341339" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 341339" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 341339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 341339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 341340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 341345" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 341345" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 341345" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 341345" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 341346" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 341403" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 341403" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 341403" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 341403" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 341404" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 342159" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 342159" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 342159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 342159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 342160" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 342160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 342181" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 342181" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 342181" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 342181" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 342182" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 342249" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 342249" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 342249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 342249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 342250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 342255" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 342255" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 342255" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 342255" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 342256" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 342313" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 342313" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 342313" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 342313" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 342314" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 343069" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 343069" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 343069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 343069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 343070" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 343070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 343091" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 343091" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 343091" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 343091" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 343092" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 343159" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 343159" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 343159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 343159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 343160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 343165" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 343165" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 343165" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 343165" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 343166" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 343223" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 343223" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 343223" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 343223" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 343224" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 343979" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 343979" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 343979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 343979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 343980" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 343980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 344001" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 344001" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 344001" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 344001" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 344002" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 344069" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 344069" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 344069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 344069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 344070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 344075" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 344075" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 344075" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 344075" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 344076" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 344133" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 344133" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 344133" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 344133" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 344134" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 344889" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 344889" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 344889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 344889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 344890" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 344890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 344911" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 344911" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 344911" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 344911" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 344912" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 344979" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 344979" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 344979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 344979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 344980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 344985" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 344985" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 344985" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 344985" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 344986" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 345043" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 345043" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 345043" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 345043" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 345044" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 345799" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 345799" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 345799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 345799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 345800" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 345800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 345821" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 345821" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 345821" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 345821" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 345822" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 345889" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 345889" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 345889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 345889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 345890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 345895" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 345895" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 345895" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 345895" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 345896" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 345953" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 345953" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 345953" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 345953" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 345954" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 346709" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 346709" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 346709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 346709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 346710" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 346710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 346731" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 346731" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 346731" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 346731" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 346732" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 346799" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 346799" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 346799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 346799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 346800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 346805" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 346805" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 346805" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 346805" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 346806" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 346863" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 346863" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 346863" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 346863" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 346864" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 347619" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 347619" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 347619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 347619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 347620" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 347620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 347641" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 347641" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 347641" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 347641" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 347642" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 347709" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 347709" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 347709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 347709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 347710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 347715" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 347715" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 347715" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 347715" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 347716" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 347773" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 347773" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 347773" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 347773" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 347774" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 348529" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 348529" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 348529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 348529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 348530" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 348530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 348551" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 348551" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 348551" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 348551" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 348552" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 348619" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 348619" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 348619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 348619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 348620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 348625" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 348625" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 348625" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 348625" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 348626" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 348683" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 348683" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 348683" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 348683" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 348684" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 349439" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 349439" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 349439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 349439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 349440" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 349440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 349461" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 349461" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 349461" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 349461" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 349462" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 349529" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 349529" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 349529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 349529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 349530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 349535" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 349535" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 349535" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 349535" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 349536" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 349593" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 349593" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 349593" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 349593" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 349594" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 350349" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 350349" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 350349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 350349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 350350" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 350350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 350371" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 350371" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 350371" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 350371" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 350372" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 350439" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 350439" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 350439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 350439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 350440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 350445" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 350445" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 350445" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 350445" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 350446" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 350503" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 350503" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 350503" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 350503" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 350504" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 351259" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 351259" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 351259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 351259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 351260" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 351260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 351281" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 351281" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 351281" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 351281" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 351282" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 351349" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 351349" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 351349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 351349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 351350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 351355" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 351355" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 351355" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 351355" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 351356" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 351413" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 351413" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 351413" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 351413" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 351414" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 352169" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 352169" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 352169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 352169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 352170" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 352170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 352191" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 352191" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 352191" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 352191" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 352192" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 352259" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 352259" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 352259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 352259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 352260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 352265" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 352265" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 352265" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 352265" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 352266" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 352323" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 352323" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 352323" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 352323" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 352324" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 353079" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 353079" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 353079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 353079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 353080" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 353080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 353101" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 353101" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 353101" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 353101" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 353102" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 353169" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 353169" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 353169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 353169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 353170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 353175" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 353175" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 353175" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 353175" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 353176" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 353233" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 353233" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 353233" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 353233" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 353234" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 353989" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 353989" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 353989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 353989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 353990" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 353990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 354011" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 354011" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 354011" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 354011" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 354012" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 354079" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 354079" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 354079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 354079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 354080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 354085" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 354085" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 354085" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 354085" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 354086" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 354143" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 354143" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 354143" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 354143" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 354144" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 354899" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 354899" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 354899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 354899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 354900" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 354900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 354921" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 354921" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 354921" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 354921" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 354922" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 354989" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 354989" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 354989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 354989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 354990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 354995" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 354995" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 354995" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 354995" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 354996" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 355053" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 355053" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 355053" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 355053" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 355054" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 355809" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 355809" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 355809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 355809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 355810" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 355810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 355831" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 355831" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 355831" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 355831" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 355832" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 355899" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 355899" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 355899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 355899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 355900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 355905" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 355905" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 355905" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 355905" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 355906" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 355963" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 355963" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 355963" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 355963" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 355964" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 356719" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 356719" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 356719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 356719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 356720" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 356720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 356741" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 356741" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 356741" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 356741" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 356742" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 356809" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 356809" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 356809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 356809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 356810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 356815" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 356815" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 356815" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 356815" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 356816" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 356873" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 356873" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 356873" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 356873" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 356874" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 357629" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 357629" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 357629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 357629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 357630" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 357630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 357651" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 357651" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 357651" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 357651" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 357652" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 357719" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 357719" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 357719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 357719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 357720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 357725" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 357725" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 357725" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 357725" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 357726" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 357783" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 357783" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 357783" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 357783" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 357784" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 358539" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 358539" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 358539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 358539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 358540" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 358540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 358561" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 358561" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 358561" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 358561" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 358562" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 358629" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 358629" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 358629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 358629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 358630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 358635" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 358635" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 358635" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 358635" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 358636" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 358693" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 358693" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 358693" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 358693" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 358694" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 359449" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 359449" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 359449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 359449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 359450" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 359450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 359471" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 359471" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 359471" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 359471" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 359472" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 359539" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 359539" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 359539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 359539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 359540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 359545" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 359545" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 359545" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 359545" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 359546" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 359603" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 359603" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 359603" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 359603" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 359604" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 360359" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 360359" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 360359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 360359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 360360" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 360360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 360381" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 360381" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 360381" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 360381" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 360382" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 360449" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 360449" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 360449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 360449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 360450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 360455" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 360455" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 360455" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 360455" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 360456" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 360513" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 360513" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 360513" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 360513" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 360514" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 361269" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 361269" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 361269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 361269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 361270" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 361270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 361291" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 361291" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 361291" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 361291" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 361292" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 361359" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 361359" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 361359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 361359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 361360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 361365" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 361365" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 361365" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 361365" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 361366" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 361423" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 361423" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 361423" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 361423" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 361424" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 362179" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 362179" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 362179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 362179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 362180" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 362180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 362201" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 362201" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 362201" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 362201" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 362202" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 362269" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 362269" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 362269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 362269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 362270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 362275" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 362275" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 362275" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 362275" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 362276" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 362333" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 362333" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 362333" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 362333" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 362334" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 363089" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 363089" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 363089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 363089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 363090" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 363090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 363111" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 363111" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 363111" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 363111" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 363112" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 363179" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 363179" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 363179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 363179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 363180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 363185" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 363185" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 363185" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 363185" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 363186" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 363243" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 363243" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 363243" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 363243" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 363244" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 363999" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 363999" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 363999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 363999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 364000" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 364000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 364021" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 364021" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 364021" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 364021" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 364022" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 364089" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 364089" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 364089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 364089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 364090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 364095" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 364095" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 364095" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 364095" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 364096" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 364153" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 364153" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 364153" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 364153" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 364154" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 364909" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 364909" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 364909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 364909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 364910" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 364910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 364931" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 364931" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 364931" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 364931" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 364932" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 364999" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 364999" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 364999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 364999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 365000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 365005" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 365005" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 365005" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 365005" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 365006" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 365063" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 365063" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 365063" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 365063" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 365064" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 365819" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 365819" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 365819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 365819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 365820" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 365820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 365841" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 365841" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 365841" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 365841" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 365842" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 365909" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 365909" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 365909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 365909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 365910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 365915" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 365915" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 365915" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 365915" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 365916" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 365973" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 365973" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 365973" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 365973" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 365974" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 366729" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 366729" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 366729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 366729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 366730" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 366730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 366751" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 366751" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 366751" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 366751" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 366752" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 366819" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 366819" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 366819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 366819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 366820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 366825" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 366825" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 366825" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 366825" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 366826" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 366883" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 366883" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 366883" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 366883" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 366884" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 367639" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 367639" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 367639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 367639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 367640" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 367640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 367661" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 367661" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 367661" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 367661" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 367662" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 367729" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 367729" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 367729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 367729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 367730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 367735" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 367735" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 367735" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 367735" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 367736" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 367793" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 367793" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 367793" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 367793" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 367794" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 368549" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 368549" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 368549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 368549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 368550" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 368550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 368571" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 368571" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 368571" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 368571" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 368572" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 368639" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 368639" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 368639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 368639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 368640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 368645" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 368645" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 368645" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 368645" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 368646" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 368703" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 368703" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 368703" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 368703" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 368704" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 369459" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 369459" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 369459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 369459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 369460" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 369460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 369481" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 369481" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 369481" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 369481" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 369482" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 369549" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 369549" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 369549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 369549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 369550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 369555" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 369555" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 369555" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 369555" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 369556" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 369613" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 369613" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 369613" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 369613" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 369614" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 370369" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 370369" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 370369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 370369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 370370" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 370370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 370391" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 370391" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 370391" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 370391" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 370392" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 370459" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 370459" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 370459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 370459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 370460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 370465" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 370465" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 370465" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 370465" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 370466" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 370523" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 370523" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 370523" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 370523" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 370524" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 371279" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 371279" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 371279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 371279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 371280" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 371280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 371301" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 371301" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 371301" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 371301" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 371302" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 371369" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 371369" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 371369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 371369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 371370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 371375" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 371375" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 371375" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 371375" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 371376" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 371433" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 371433" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 371433" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 371433" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 371434" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 372189" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 372189" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 372189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 372189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 372190" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 372190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 372211" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 372211" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 372211" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 372211" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 372212" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 372279" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 372279" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 372279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 372279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 372280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 372285" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 372285" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 372285" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 372285" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 372286" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 372343" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 372343" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 372343" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 372343" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 372344" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 373099" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 373099" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 373099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 373099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 373100" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 373100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 373121" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 373121" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 373121" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 373121" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 373122" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 373189" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 373189" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 373189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 373189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 373190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 373195" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 373195" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 373195" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 373195" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 373196" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 373253" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 373253" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 373253" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 373253" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 373254" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 374009" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 374009" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 374009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 374009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 374010" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 374010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 374031" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 374031" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 374031" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 374031" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 374032" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 374099" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 374099" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 374099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 374099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 374100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 374105" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 374105" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 374105" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 374105" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 374106" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 374163" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 374163" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 374163" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 374163" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 374164" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 374919" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 374919" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 374919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 374919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 374920" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 374920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 374941" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 374941" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 374941" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 374941" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 374942" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 375009" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 375009" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 375009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 375009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 375010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 375015" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 375015" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 375015" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 375015" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 375016" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 375073" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 375073" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 375073" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 375073" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 375074" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 375829" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 375829" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 375829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 375829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 375830" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 375830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 375851" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 375851" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 375851" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 375851" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 375852" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 375919" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 375919" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 375919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 375919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 375920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 375925" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 375925" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 375925" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 375925" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 375926" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 375983" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 375983" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 375983" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 375983" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 375984" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 376739" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 376739" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 376739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 376739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 376740" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 376740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 376761" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 376761" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 376761" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 376761" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 376762" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 376829" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 376829" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 376829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 376829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 376830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 376835" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 376835" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 376835" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 376835" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 376836" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 376893" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 376893" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 376893" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 376893" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 376894" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 377649" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 377649" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 377649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 377649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 377650" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 377650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 377671" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 377671" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 377671" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 377671" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 377672" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 377739" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 377739" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 377739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 377739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 377740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 377745" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 377745" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 377745" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 377745" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 377746" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 377803" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 377803" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 377803" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 377803" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 377804" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 378559" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 378559" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 378559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 378559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 378560" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 378560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 378581" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 378581" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 378581" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 378581" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 378582" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 378649" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 378649" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 378649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 378649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 378650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 378655" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 378655" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 378655" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 378655" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 378656" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 378713" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 378713" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 378713" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 378713" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 378714" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 379469" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 379469" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 379469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 379469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 379470" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 379470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 379491" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 379491" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 379491" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 379491" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 379492" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 379559" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 379559" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 379559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 379559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 379560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 379565" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 379565" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 379565" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 379565" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 379566" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 379623" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 379623" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 379623" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 379623" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 379624" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 380379" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 380379" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 380379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 380379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 380380" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 380380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 380401" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 380401" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 380401" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 380401" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 380402" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 380469" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 380469" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 380469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 380469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 380470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 380475" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 380475" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 380475" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 380475" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 380476" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 380533" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 380533" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 380533" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 380533" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 380534" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 381289" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 381289" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 381289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 381289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 381290" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 381290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 381311" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 381311" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 381311" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 381311" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 381312" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 381379" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 381379" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 381379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 381379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 381380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 381385" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 381385" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 381385" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 381385" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 381386" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 381443" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 381443" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 381443" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 381443" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 381444" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 382199" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 382199" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 382199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 382199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 382200" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 382200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 382221" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 382221" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 382221" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 382221" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 382222" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 382289" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 382289" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 382289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 382289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 382290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 382295" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 382295" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 382295" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 382295" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 382296" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 382353" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 382353" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 382353" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 382353" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 382354" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 383109" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 383109" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 383109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 383109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 383110" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 383110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 383131" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 383131" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 383131" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 383131" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 383132" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 383199" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 383199" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 383199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 383199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 383200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 383205" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 383205" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 383205" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 383205" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 383206" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 383263" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 383263" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 383263" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 383263" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 383264" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 384019" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 384019" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 384019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 384019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 384020" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 384020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 384041" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 384041" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 384041" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 384041" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 384042" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 384109" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 384109" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 384109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 384109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 384110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 384115" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 384115" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 384115" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 384115" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 384116" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 384173" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 384173" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 384173" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 384173" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 384174" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 384929" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 384929" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 384929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 384929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 384930" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 384930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 384951" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 384951" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 384951" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 384951" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 384952" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 385019" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 385019" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 385019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 385019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 385020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 385025" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 385025" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 385025" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 385025" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 385026" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 385083" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 385083" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 385083" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 385083" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 385084" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 385839" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 385839" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 385839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 385839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 385840" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 385840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 385861" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 385861" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 385861" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 385861" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 385862" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 385929" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 385929" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 385929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 385929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 385930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 385935" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 385935" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 385935" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 385935" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 385936" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 385993" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 385993" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 385993" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 385993" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 385994" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 386749" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 386749" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 386749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 386749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 386750" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 386750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 386771" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 386771" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 386771" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 386771" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 386772" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 386839" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 386839" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 386839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 386839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 386840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 386845" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 386845" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 386845" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 386845" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 386846" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 386903" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 386903" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 386903" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 386903" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 386904" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 387659" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 387659" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 387659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 387659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 387660" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 387660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 387681" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 387681" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 387681" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 387681" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 387682" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 387749" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 387749" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 387749" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 387749" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 387750" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 387755" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 387755" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 387755" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 387755" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 387756" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 387813" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 387813" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 387813" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 387813" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 387814" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 388569" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 388569" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 388569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 388569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 388570" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 388570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 388591" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 388591" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 388591" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 388591" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 388592" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 388659" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 388659" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 388659" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 388659" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 388660" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 388665" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 388665" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 388665" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 388665" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 388666" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 388723" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 388723" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 388723" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 388723" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 388724" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 389479" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 389479" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 389479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 389479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 389480" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 389480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 389501" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 389501" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 389501" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 389501" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 389502" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 389569" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 389569" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 389569" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 389569" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 389570" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 389575" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 389575" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 389575" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 389575" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 389576" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 389633" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 389633" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 389633" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 389633" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 389634" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 390389" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 390389" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 390389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 390389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 390390" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 390390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 390411" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 390411" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 390411" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 390411" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 390412" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 390479" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 390479" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 390479" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 390479" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 390480" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 390485" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 390485" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 390485" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 390485" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 390486" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 390543" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 390543" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 390543" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 390543" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 390544" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 391299" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 391299" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 391299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 391299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 391300" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 391300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 391321" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 391321" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 391321" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 391321" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 391322" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 391389" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 391389" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 391389" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 391389" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 391390" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 391395" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 391395" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 391395" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 391395" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 391396" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 391453" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 391453" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 391453" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 391453" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 391454" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 392209" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 392209" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 392209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 392209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 392210" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 392210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 392231" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 392231" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 392231" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 392231" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 392232" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 392299" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 392299" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 392299" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 392299" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 392300" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 392305" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 392305" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 392305" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 392305" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 392306" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 392363" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 392363" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 392363" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 392363" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 392364" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 393119" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 393119" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 393119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 393119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 393120" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 393120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 393141" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 393141" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 393141" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 393141" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 393142" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 393209" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 393209" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 393209" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 393209" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 393210" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 393215" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 393215" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 393215" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 393215" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 393216" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 393273" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 393273" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 393273" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 393273" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 393274" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 394029" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 394029" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 394029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 394029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 394030" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 394030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 394051" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 394051" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 394051" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 394051" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 394052" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 394119" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 394119" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 394119" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 394119" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 394120" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 394125" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 394125" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 394125" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 394125" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 394126" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 394183" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 394183" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 394183" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 394183" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 394184" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 394939" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 394939" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 394939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 394939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 394940" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 394940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 394961" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 394961" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 394961" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 394961" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 394962" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 395029" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 395029" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 395029" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 395029" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 395030" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 395035" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 395035" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 395035" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 395035" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 395036" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 395093" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 395093" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 395093" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 395093" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 395094" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 395849" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 395849" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 395849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 395849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 395850" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 395850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 395871" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 395871" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 395871" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 395871" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 395872" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 395939" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 395939" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 395939" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 395939" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 395940" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 395945" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 395945" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 395945" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 395945" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 395946" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 396003" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 396003" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 396003" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 396003" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 396004" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 396759" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 396759" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 396759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 396759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 396760" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 396760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 396781" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 396781" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 396781" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 396781" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 396782" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 396849" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 396849" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 396849" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 396849" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 396850" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 396855" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 396855" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 396855" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 396855" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 396856" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 396913" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 396913" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 396913" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 396913" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 396914" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 397669" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 397669" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 397669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 397669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 397670" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 397670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 397691" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 397691" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 397691" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 397691" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 397692" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 397759" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 397759" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 397759" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 397759" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 397760" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 397765" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 397765" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 397765" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 397765" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 397766" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 397823" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 397823" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 397823" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 397823" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 397824" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 398579" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 398579" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 398579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 398579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 398580" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 398580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 398601" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 398601" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 398601" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 398601" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 398602" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 398669" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 398669" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 398669" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 398669" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 398670" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 398675" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 398675" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 398675" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 398675" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 398676" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 398733" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 398733" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 398733" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 398733" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 398734" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 399489" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 399489" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 399489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 399489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 399490" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 399490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 399511" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 399511" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 399511" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 399511" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 399512" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 399579" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 399579" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 399579" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 399579" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 399580" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 399585" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 399585" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 399585" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 399585" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 399586" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 399643" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 399643" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 399643" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 399643" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 399644" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 400399" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 400399" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 400399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 400399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 400400" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 400400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 400421" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 400421" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 400421" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 400421" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 400422" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 400489" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 400489" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 400489" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 400489" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 400490" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 400495" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 400495" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 400495" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 400495" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 400496" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 400553" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 400553" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 400553" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 400553" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 400554" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 401309" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 401309" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 401309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 401309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 401310" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 401310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 401331" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 401331" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 401331" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 401331" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 401332" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 401399" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 401399" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 401399" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 401399" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 401400" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 401405" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 401405" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 401405" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 401405" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 401406" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 401463" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 401463" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 401463" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 401463" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 401464" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 402219" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 402219" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 402219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 402219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 402220" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 402220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 402241" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 402241" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 402241" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 402241" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 402242" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 402309" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 402309" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 402309" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 402309" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 402310" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 402315" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 402315" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 402315" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 402315" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 402316" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 402373" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 402373" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 402373" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 402373" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 402374" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 403129" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 403129" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 403129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 403129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 403130" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 403130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 403151" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 403151" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 403151" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 403151" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 403152" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 403219" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 403219" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 403219" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 403219" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 403220" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 403225" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 403225" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 403225" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 403225" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 403226" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 403283" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 403283" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 403283" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 403283" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 403284" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 404039" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 404039" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 404039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 404039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 404040" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 404040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 404061" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 404061" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 404061" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 404061" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 404062" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 404129" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 404129" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 404129" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 404129" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 404130" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 404135" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 404135" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 404135" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 404135" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 404136" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 404193" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 404193" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 404193" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 404193" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 404194" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 404949" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 404949" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 404949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 404949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 404950" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 404950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 404971" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 404971" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 404971" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 404971" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 404972" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 405039" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 405039" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 405039" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 405039" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 405040" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 405045" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 405045" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 405045" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 405045" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 405046" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 405103" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 405103" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 405103" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 405103" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 405104" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 405859" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 405859" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 405859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 405859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 405860" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 405860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 405881" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 405881" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 405881" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 405881" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 405882" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 405949" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 405949" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 405949" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 405949" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 405950" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 405955" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 405955" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 405955" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 405955" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 405956" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 406013" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 406013" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 406013" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 406013" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 406014" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 406769" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 406769" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 406769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 406769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 406770" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 406770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 406791" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 406791" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 406791" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 406791" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 406792" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 406859" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 406859" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 406859" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 406859" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 406860" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 406865" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 406865" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 406865" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 406865" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 406866" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 406923" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 406923" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 406923" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 406923" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 406924" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 407679" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 407679" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 407679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 407679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 407680" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 407680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 407701" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 407701" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 407701" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 407701" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 407702" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 407769" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 407769" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 407769" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 407769" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 407770" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 407775" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 407775" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 407775" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 407775" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 407776" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 407833" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 407833" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 407833" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 407833" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 407834" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 408589" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 408589" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 408589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 408589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 408590" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 408590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 408611" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 408611" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 408611" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 408611" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 408612" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 408679" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 408679" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 408679" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 408679" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 408680" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 408685" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 408685" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 408685" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 408685" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 408686" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 408743" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 408743" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 408743" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 408743" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 408744" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 409499" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 409499" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 409499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 409499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 409500" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 409500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 409521" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 409521" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 409521" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 409521" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 409522" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 409589" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 409589" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 409589" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 409589" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 409590" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 409595" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 409595" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 409595" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 409595" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 409596" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 409653" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 409653" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 409653" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 409653" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 409654" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 410409" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 410409" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 410409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 410409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 410410" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 410410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 410431" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 410431" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 410431" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 410431" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 410432" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 410499" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 410499" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 410499" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 410499" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 410500" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 410505" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 410505" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 410505" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 410505" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 410506" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 410563" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 410563" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 410563" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 410563" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 410564" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 411319" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 411319" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 411319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 411319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 411320" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 411320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 411341" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 411341" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 411341" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 411341" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 411342" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 411409" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 411409" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 411409" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 411409" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 411410" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 411415" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 411415" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 411415" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 411415" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 411416" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 411473" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 411473" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 411473" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 411473" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 411474" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 412229" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 412229" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 412229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 412229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 412230" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 412230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 412251" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 412251" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 412251" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 412251" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 412252" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 412319" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 412319" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 412319" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 412319" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 412320" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 412325" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 412325" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 412325" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 412325" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 412326" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 412383" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 412383" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 412383" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 412383" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 412384" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 413139" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 413139" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 413139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 413139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 413140" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 413140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 413161" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 413161" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 413161" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 413161" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 413162" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 413229" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 413229" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 413229" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 413229" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 413230" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 413235" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 413235" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 413235" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 413235" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 413236" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 413293" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 413293" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 413293" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 413293" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 413294" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 414049" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 414049" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 414049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 414049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 414050" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 414050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 414071" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 414071" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 414071" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 414071" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 414072" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 414139" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 414139" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 414139" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 414139" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 414140" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 414145" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 414145" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 414145" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 414145" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 414146" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 414203" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 414203" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 414203" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 414203" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 414204" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 414959" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 414959" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 414959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 414959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 414960" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 414960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 414981" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 414981" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 414981" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 414981" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 414982" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 415049" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 415049" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 415049" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 415049" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 415050" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 415055" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 415055" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 415055" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 415055" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 415056" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 415113" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 415113" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 415113" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 415113" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 415114" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 415869" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 415869" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 415869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 415869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 415870" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 415870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 415891" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 415891" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 415891" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 415891" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 415892" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 415959" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 415959" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 415959" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 415959" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 415960" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 415965" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 415965" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 415965" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 415965" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 415966" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 416023" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 416023" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 416023" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 416023" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 416024" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 416779" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 416779" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 416779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 416779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 416780" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 416780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 416801" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 416801" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 416801" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 416801" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 416802" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 416869" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 416869" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 416869" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 416869" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 416870" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 416875" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 416875" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 416875" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 416875" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 416876" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 416933" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 416933" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 416933" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 416933" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 416934" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 417689" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 417689" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 417689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 417689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 417690" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 417690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 417711" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 417711" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 417711" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 417711" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 417712" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 417779" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 417779" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 417779" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 417779" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 417780" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 417785" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 417785" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 417785" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 417785" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 417786" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 417843" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 417843" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 417843" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 417843" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 417844" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 418599" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 418599" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 418599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 418599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 418600" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 418600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 418621" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 418621" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 418621" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 418621" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 418622" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 418689" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 418689" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 418689" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 418689" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 418690" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 418695" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 418695" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 418695" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 418695" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 418696" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 418753" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 418753" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 418753" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 418753" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 418754" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 419509" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 419509" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 419509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 419509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 419510" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 419510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 419531" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 419531" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 419531" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 419531" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 419532" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 419599" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 419599" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 419599" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 419599" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 419600" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 419605" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 419605" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 419605" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 419605" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 419606" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 419663" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 419663" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 419663" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 419663" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 419664" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 420419" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 420419" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 420419" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 420419" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 420420" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 420420" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 420441" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 420441" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 420441" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 420441" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 420442" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 420509" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 420509" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 420509" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 420509" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 420510" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 420515" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 420515" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 420515" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 420515" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 420516" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 420573" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 420573" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 420573" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 420573" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 420574" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 421329" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 421329" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 421329" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 421329" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 421330" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 421330" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 421351" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 421351" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 421351" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 421351" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 421352" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 421419" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 421419" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 421419" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 421419" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 421420" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 421425" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 421425" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 421425" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 421425" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 421426" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 421483" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 421483" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 421483" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 421483" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 421484" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 422239" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 422239" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 422239" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 422239" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 422240" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 422240" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 422261" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 422261" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 422261" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 422261" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 422262" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 422329" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 422329" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 422329" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 422329" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 422330" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 422335" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 422335" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 422335" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 422335" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 422336" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 422393" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 422393" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 422393" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 422393" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 422394" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 423149" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 423149" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 423149" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 423149" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 423150" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 423150" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 423171" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 423171" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 423171" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 423171" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 423172" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 423239" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 423239" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 423239" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 423239" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 423240" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 423245" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 423245" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 423245" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 423245" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 423246" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 423303" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 423303" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 423303" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 423303" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 423304" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 424059" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 424059" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 424059" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 424059" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 424060" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 424060" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 424081" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 424081" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 424081" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 424081" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 424082" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 424149" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 424149" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 424149" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 424149" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 424150" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 424155" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 424155" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 424155" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 424155" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 424156" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 424213" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 424213" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 424213" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 424213" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 424214" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 424969" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 424969" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 424969" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 424969" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 424970" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 424970" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 424991" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 424991" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 424991" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 424991" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 424992" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 425059" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 425059" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 425059" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 425059" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 425060" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 425065" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 425065" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 425065" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 425065" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 425066" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 425123" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 425123" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 425123" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 425123" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 425124" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 425879" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 425879" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 425879" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 425879" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 425880" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 425880" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 425901" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 425901" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 425901" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 425901" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 425902" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 425969" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 425969" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 425969" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 425969" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 425970" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 425975" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 425975" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 425975" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 425975" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 425976" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 426033" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 426033" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 426033" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 426033" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 426034" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 426789" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 426789" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 426789" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 426789" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 426790" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 426790" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 426811" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 426811" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 426811" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 426811" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 426812" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 426879" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 426879" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 426879" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 426879" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 426880" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 426885" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 426885" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 426885" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 426885" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 426886" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 426943" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 426943" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 426943" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 426943" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 426944" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 427699" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 427699" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 427699" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 427699" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 427700" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 427700" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 427721" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 427721" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 427721" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 427721" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 427722" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 427789" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 427789" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 427789" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 427789" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 427790" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 427795" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 427795" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 427795" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 427795" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 427796" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 427853" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 427853" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 427853" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 427853" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 427854" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 428609" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 428609" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 428609" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 428609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 428610" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 428610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 428631" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 428631" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 428631" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 428631" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 428632" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 428699" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 428699" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 428699" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 428699" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 428700" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 428705" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 428705" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 428705" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 428705" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 428706" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 428763" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 428763" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 428763" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 428763" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 428764" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 429519" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 429519" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 429519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 429519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 429520" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 429520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 429541" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 429541" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 429541" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 429541" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 429542" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 429609" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 429609" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 429609" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 429609" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 429610" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 429615" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 429615" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 429615" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 429615" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 429616" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 429673" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 429673" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 429673" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 429673" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 429674" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 430429" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 430429" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 430429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 430429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 430430" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 430430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 430451" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 430451" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 430451" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 430451" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 430452" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 430519" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 430519" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 430519" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 430519" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 430520" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 430525" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 430525" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 430525" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 430525" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 430526" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 430583" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 430583" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 430583" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 430583" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 430584" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 431339" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 431339" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 431339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 431339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 431340" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 431340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 431361" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 431361" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 431361" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 431361" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 431362" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 431429" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 431429" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 431429" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 431429" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 431430" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 431435" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 431435" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 431435" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 431435" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 431436" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 431493" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 431493" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 431493" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 431493" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 431494" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 432249" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 432249" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 432249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 432249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 432250" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 432250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 432271" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 432271" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 432271" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 432271" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 432272" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 432339" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 432339" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 432339" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 432339" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 432340" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 432345" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 432345" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 432345" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 432345" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 432346" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 432403" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 432403" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 432403" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 432403" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 432404" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 433159" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 433159" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 433159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 433159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 433160" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 433160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 433181" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 433181" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 433181" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 433181" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 433182" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 433249" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 433249" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 433249" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 433249" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 433250" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 433255" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 433255" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 433255" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 433255" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 433256" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 433313" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 433313" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 433313" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 433313" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 433314" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 434069" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 434069" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 434069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 434069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 434070" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 434070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 434091" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 434091" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 434091" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 434091" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 434092" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 434159" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 434159" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 434159" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 434159" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 434160" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 434165" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 434165" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 434165" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 434165" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 434166" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 434223" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 434223" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 434223" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 434223" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 434224" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 434979" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 434979" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 434979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 434979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 434980" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 434980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 435001" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 435001" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 435001" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 435001" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 435002" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 435069" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 435069" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 435069" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 435069" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 435070" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 435075" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 435075" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 435075" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 435075" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 435076" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 435133" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 435133" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 435133" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 435133" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 435134" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 435889" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 435889" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 435889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 435889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 435890" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 435890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 435911" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 435911" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 435911" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 435911" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 435912" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 435979" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 435979" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 435979" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 435979" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 435980" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 435985" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 435985" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 435985" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 435985" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 435986" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 436043" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 436043" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 436043" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 436043" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 436044" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 436799" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 436799" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 436799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 436799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 436800" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 436800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 436821" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 436821" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 436821" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 436821" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 436822" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 436889" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 436889" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 436889" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 436889" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 436890" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 436895" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 436895" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 436895" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 436895" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 436896" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 436953" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 436953" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 436953" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 436953" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 436954" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 437709" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 437709" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 437709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 437709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 437710" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 437710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 437731" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 437731" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 437731" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 437731" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 437732" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 437799" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 437799" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 437799" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 437799" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 437800" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 437805" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 437805" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 437805" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 437805" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 437806" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 437863" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 437863" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 437863" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 437863" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 437864" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 438619" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 438619" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 438619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 438619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 438620" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 438620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 438641" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 438641" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 438641" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 438641" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 438642" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 438709" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 438709" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 438709" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 438709" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 438710" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 438715" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 438715" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 438715" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 438715" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 438716" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 438773" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 438773" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 438773" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 438773" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 438774" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 439529" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 439529" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 439529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 439529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 439530" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 439530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 439551" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 439551" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 439551" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 439551" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 439552" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 439619" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 439619" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 439619" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 439619" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 439620" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 439625" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 439625" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 439625" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 439625" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 439626" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 439683" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 439683" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 439683" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 439683" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 439684" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 440439" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 440439" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 440439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 440439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 440440" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 440440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 440461" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 440461" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 440461" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 440461" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 440462" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 440529" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 440529" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 440529" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 440529" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 440530" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 440535" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 440535" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 440535" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 440535" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 440536" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 440593" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 440593" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 440593" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 440593" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 440594" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 441349" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 441349" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 441349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 441349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 441350" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 441350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 441371" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 441371" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 441371" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 441371" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 441372" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 441439" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 441439" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 441439" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 441439" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 441440" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 441445" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 441445" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 441445" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 441445" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 441446" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 441503" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 441503" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 441503" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 441503" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 441504" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 442259" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 442259" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 442259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 442259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 442260" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 442260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 442281" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 442281" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 442281" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 442281" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 442282" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 442349" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 442349" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 442349" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 442349" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 442350" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 442355" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 442355" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 442355" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 442355" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 442356" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 442413" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 442413" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 442413" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 442413" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 442414" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 443169" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 443169" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 443169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 443169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 443170" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 443170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 443191" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 443191" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 443191" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 443191" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 443192" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 443259" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 443259" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 443259" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 443259" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 443260" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 443265" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 443265" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 443265" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 443265" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 443266" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 443323" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 443323" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 443323" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 443323" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 443324" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 444079" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 444079" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 444079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 444079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 444080" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 444080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 444101" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 444101" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 444101" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 444101" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 444102" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 444169" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 444169" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 444169" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 444169" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 444170" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 444175" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 444175" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 444175" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 444175" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 444176" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 444233" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 444233" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 444233" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 444233" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 444234" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 444989" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 444989" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 444989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 444989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 444990" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 444990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 445011" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 445011" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 445011" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 445011" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 445012" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 445079" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 445079" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 445079" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 445079" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 445080" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 445085" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 445085" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 445085" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 445085" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 445086" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 445143" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 445143" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 445143" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 445143" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 445144" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 445899" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 445899" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 445899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 445899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 445900" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 445900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 445921" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 445921" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 445921" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 445921" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 445922" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 445989" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 445989" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 445989" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 445989" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 445990" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 445995" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 445995" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 445995" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 445995" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 445996" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 446053" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 446053" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 446053" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 446053" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 446054" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 446809" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 446809" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 446809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 446809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 446810" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 446810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 446831" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 446831" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 446831" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 446831" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 446832" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 446899" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 446899" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 446899" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 446899" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 446900" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 446905" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 446905" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 446905" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 446905" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 446906" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 446963" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 446963" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 446963" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 446963" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 446964" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 447719" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 447719" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 447719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 447719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 447720" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 447720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 447741" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 447741" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 447741" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 447741" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 447742" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 447809" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 447809" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 447809" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 447809" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 447810" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 447815" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 447815" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 447815" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 447815" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 447816" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 447873" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 447873" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 447873" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 447873" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 447874" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 448629" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 448629" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 448629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 448629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 448630" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 448630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 448651" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 448651" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 448651" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 448651" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 448652" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 448719" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 448719" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 448719" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 448719" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 448720" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 448725" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 448725" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 448725" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 448725" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 448726" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 448783" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 448783" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 448783" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 448783" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 448784" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 449539" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 449539" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 449539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 449539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 449540" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 449540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 449561" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 449561" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 449561" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 449561" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 449562" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 449629" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 449629" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 449629" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 449629" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 449630" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 449635" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 449635" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 449635" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 449635" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 449636" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 449693" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 449693" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 449693" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 449693" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 449694" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 450449" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 450449" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 450449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 450449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 450450" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 450450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 450471" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 450471" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 450471" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 450471" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 450472" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 450539" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 450539" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 450539" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 450539" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 450540" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 450545" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 450545" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 450545" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 450545" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 450546" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 450603" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 450603" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 450603" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 450603" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 450604" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 451359" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 451359" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 451359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 451359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 451360" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 451360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 451381" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 451381" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 451381" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 451381" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 451382" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 451449" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 451449" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 451449" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 451449" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 451450" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 451455" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 451455" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 451455" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 451455" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 451456" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 451513" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 451513" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 451513" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 451513" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 451514" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 452269" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 452269" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 452269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 452269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 452270" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 452270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 452291" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 452291" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 452291" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 452291" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 452292" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 452359" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 452359" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 452359" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 452359" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 452360" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 452365" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 452365" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 452365" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 452365" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 452366" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 452423" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 452423" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 452423" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 452423" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 452424" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 453179" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 453179" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 453179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 453179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 453180" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 453180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 453201" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 453201" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 453201" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 453201" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 453202" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 453269" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 453269" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 453269" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 453269" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 453270" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 453275" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 453275" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 453275" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 453275" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 453276" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 453333" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 453333" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 453333" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 453333" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 453334" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 454089" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 454089" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 454089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 454089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 454090" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 454090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 454111" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 454111" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 454111" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 454111" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 454112" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 454179" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 454179" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 454179" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 454179" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 454180" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 454185" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 454185" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 454185" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 454185" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 454186" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 454243" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 454243" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 454243" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 454243" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 454244" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 454999" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 454999" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 454999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 454999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 455000" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 455000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 455021" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 455021" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 455021" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 455021" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 455022" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 455089" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 455089" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 455089" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 455089" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 455090" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 455095" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 455095" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 455095" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 455095" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 455096" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 455153" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 455153" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 455153" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 455153" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 455154" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 455909" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 455909" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 455909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 455909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 455910" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 455910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 455931" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 455931" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 455931" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 455931" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 455932" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 455999" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 455999" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 455999" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 455999" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 456000" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 456005" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 456005" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 456005" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 456005" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 456006" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 456063" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 456063" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 456063" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 456063" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 456064" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 456819" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 456819" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 456819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 456819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 456820" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 456820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 456841" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 456841" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 456841" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 456841" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 456842" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 456909" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 456909" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 456909" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 456909" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 456910" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 456915" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 456915" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 456915" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 456915" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 456916" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 456973" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 456973" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 456973" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 456973" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 456974" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 457729" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 457729" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 457729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 457729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 457730" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 457730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 457751" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 457751" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 457751" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 457751" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 457752" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 457819" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 457819" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 457819" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 457819" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 457820" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 457825" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 457825" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 457825" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 457825" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 457826" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 457883" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 457883" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 457883" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 457883" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 457884" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 458639" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 458639" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 458639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 458639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 458640" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 458640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 458661" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 458661" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 458661" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 458661" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 458662" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 458729" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 458729" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 458729" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 458729" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 458730" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 458735" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 458735" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 458735" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 458735" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 458736" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 458793" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 458793" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 458793" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 458793" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 458794" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 459549" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 459549" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 459549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 459549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 459550" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 459550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 459571" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 459571" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 459571" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 459571" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 459572" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 459639" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 459639" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 459639" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 459639" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 459640" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 459645" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 459645" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 459645" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 459645" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 459646" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 459703" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 459703" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 459703" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 459703" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 459704" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 460459" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 460459" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 460459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 460459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 460460" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 460460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 460481" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 460481" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 460481" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 460481" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 460482" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 460549" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 460549" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 460549" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 460549" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 460550" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 460555" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 460555" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 460555" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 460555" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 460556" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 460613" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 460613" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 460613" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 460613" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 460614" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 461369" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 461369" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 461369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 461369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 461370" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 461370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 461391" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 461391" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 461391" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 461391" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 461392" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 461459" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 461459" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 461459" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 461459" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 461460" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 461465" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 461465" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 461465" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 461465" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 461466" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 461523" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 461523" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 461523" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 461523" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 461524" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 462279" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 462279" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 462279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 462279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 462280" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 462280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 462301" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 462301" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 462301" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 462301" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 462302" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 462369" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 462369" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 462369" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 462369" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 462370" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 462375" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 462375" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 462375" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 462375" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 462376" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 462433" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 462433" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 462433" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 462433" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 462434" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 463189" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 463189" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 463189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 463189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 463190" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 463190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 463211" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 463211" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 463211" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 463211" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 463212" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 463279" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 463279" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 463279" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 463279" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 463280" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 463285" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 463285" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 463285" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 463285" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 463286" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 463343" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 463343" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 463343" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 463343" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 463344" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 464099" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 464099" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 464099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 464099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 464100" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 464100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 464121" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 464121" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 464121" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 464121" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 464122" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 464189" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 464189" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 464189" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 464189" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 464190" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 464195" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 464195" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 464195" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 464195" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 464196" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 464253" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 464253" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 464253" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 464253" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 464254" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 465009" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 465009" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 465009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 465009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 465010" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 465010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 465031" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 465031" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 465031" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 465031" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 465032" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 465099" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 465099" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 465099" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 465099" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 465100" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 465105" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 465105" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 465105" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 465105" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 465106" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 465163" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 465163" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 465163" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 465163" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 465164" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 465919" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 465919" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 465919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 465919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 465920" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 465920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 465941" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 465941" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 465941" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 465941" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 465942" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 466009" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 466009" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 466009" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 466009" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 466010" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 466015" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 466015" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 466015" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 466015" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 466016" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 466073" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 466073" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 466073" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 466073" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 466074" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 466829" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 466829" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 466829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 466829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 466830" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 466830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 466851" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 466851" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 466851" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 466851" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 466852" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 466919" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 466919" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 466919" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 466919" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 466920" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 466925" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 466925" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 466925" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 466925" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 466926" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 466983" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 466983" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 466983" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 466983" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 466984" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 467739" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 467739" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 467739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 467739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 467740" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 467740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 467761" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 467761" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 467761" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 467761" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 467762" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 467829" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 467829" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 467829" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 467829" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 467830" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 467835" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 467835" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 467835" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 467835" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 467836" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 467893" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 467893" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 467893" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 467893" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 467894" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 468649" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 468649" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 468649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 468649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 468650" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 468650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 468671" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 468671" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 468671" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 468671" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 468672" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 468739" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 468739" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 468739" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 468739" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 468740" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 468745" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 468745" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 468745" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 468745" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 468746" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 468803" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 468803" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 468803" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 468803" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 468804" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 469559" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 469559" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 469559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 469559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 469560" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 469560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 469581" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 469581" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 469581" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 469581" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 469582" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 469649" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 469649" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 469649" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 469649" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 469650" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 469655" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 469655" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 469655" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 469655" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 469656" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 469713" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 469713" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 469713" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 469713" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 469714" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 470469" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 470469" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 470469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 470469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 470470" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 470470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 470491" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 470491" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 470491" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 470491" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 470492" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 470559" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 470559" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 470559" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 470559" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 470560" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 470565" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 470565" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 470565" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 470565" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 470566" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 470623" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 470623" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 470623" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 470623" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 470624" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 471379" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 471379" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 471379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 471379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 471380" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 471380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 471401" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 471401" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 471401" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 471401" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 471402" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 471469" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 471469" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 471469" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 471469" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 471470" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 471475" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 471475" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 471475" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 471475" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 471476" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 471533" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 471533" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 471533" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 471533" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 471534" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 472289" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 472289" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 472289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 472289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 472290" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 472290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 472311" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 472311" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 472311" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 472311" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 472312" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 472379" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 472379" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 472379" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 472379" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 472380" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 472385" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 472385" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 472385" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 472385" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 472386" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 472443" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 472443" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 472443" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 472443" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 472444" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 473199" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 473199" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 473199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 473199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 473200" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 473200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 473221" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 473221" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 473221" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 473221" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 473222" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 473289" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 473289" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 473289" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 473289" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 473290" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 473295" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 473295" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 473295" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 473295" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 473296" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 473353" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 473353" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 473353" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 473353" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 473354" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 474109" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 474109" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 474109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 474109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 474110" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 474110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 474131" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 474131" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 474131" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 474131" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 474132" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 474199" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 474199" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 474199" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 474199" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 474200" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 474205" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 474205" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 474205" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 474205" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 474206" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 474263" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 474263" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 474263" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 474263" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 474264" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 475019" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 475019" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 475019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 475019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 475020" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 475020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 475041" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 475041" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 475041" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 475041" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 475042" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 475109" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 475109" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 475109" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 475109" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 475110" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 475115" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 475115" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 475115" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 475115" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 475116" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 475173" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 475173" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 475173" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 475173" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 475174" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 475929" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 475929" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 475929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 475929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 475930" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 475930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 475951" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 475951" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 475951" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 475951" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 475952" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 476019" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 476019" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 476019" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 476019" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 476020" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 476025" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 476025" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 476025" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 476025" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 476026" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 476083" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 476083" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 476083" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 476083" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 476084" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 755);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 476839" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 476839" severity error;
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 476839" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 476839" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 476840" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 476840" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 21);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 476861" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 476861" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 476861" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 476861" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 476862" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 67);
		assert (csync_prime = '0') report "Unexpected value for csync_prime at cycle 476929" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 476929" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 476929" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 476929" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 476930" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 5);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 476935" severity error;
		assert (hsync2_prime = '0') report "Unexpected value for hsync2_prime at cycle 476935" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 476935" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 476935" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 476936" severity error;

		--making sure existing signals haven't changed prematurely
		wait for (clock14_3_period * 57);
		assert (csync_prime = '1') report "Unexpected value for csync_prime at cycle 476993" severity error;
		assert (hsync2_prime = '1') report "Unexpected value for hsync2_prime at cycle 476993" severity error;
		assert (sgblk_prime = '0') report "Unexpected value for sgblk_prime at cycle 476993" severity error;
		assert (vsync2_prime = '1') report "Unexpected value for vsync2_prime at cycle 476993" severity error;
		wait for clock14_3_period;

		--next cycle transition
		assert (sgblk_prime = '1') report "Unexpected value for sgblk_prime at cycle 476994" severity error;

      wait;
   end process;

END;
